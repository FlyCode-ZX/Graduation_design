always@(posedge CLK)begin


BRAM[0]<= 32'h2000A080;
BRAM[1]<= 32'h000000ED;
BRAM[2]<= 32'h000000F5;
BRAM[3]<= 32'h000000FD;
BRAM[4]<= 32'h00000105;
BRAM[5]<= 32'h0000010D;
BRAM[6]<= 32'h00000115;
BRAM[7]<= 32'h00000000;
BRAM[8]<= 32'h00000000;
BRAM[9]<= 32'h00000000;
BRAM[10]<= 32'h00000000;
BRAM[11]<= 32'h0000011D;
BRAM[12]<= 32'h00000125;
BRAM[13]<= 32'h00000000;
BRAM[14]<= 32'h0000012D;
BRAM[15]<= 32'h00000135;
BRAM[16]<= 32'h0000013D;
BRAM[17]<= 32'h00000145;
BRAM[18]<= 32'h0000014D;
BRAM[19]<= 32'h00000155;
BRAM[20]<= 32'hF802F000;
BRAM[21]<= 32'hF83AF000;
BRAM[22]<= 32'hE890A00A;
BRAM[23]<= 32'h44820C00;
BRAM[24]<= 32'hF1AA4483;
BRAM[25]<= 32'h45DA0701;
BRAM[26]<= 32'hF000D101;
BRAM[27]<= 32'hF2AFF82F;
BRAM[28]<= 32'hE8BA0E09;
BRAM[29]<= 32'hF013000F;
BRAM[30]<= 32'hBF180F01;
BRAM[31]<= 32'hF0431AFB;
BRAM[32]<= 32'h47180301;
BRAM[33]<= 32'h000046F4;
BRAM[34]<= 32'h00004714;
BRAM[35]<= 32'hBF243A10;
BRAM[36]<= 32'hC178C878;
BRAM[37]<= 32'h0752D8FA;
BRAM[38]<= 32'hC830BF24;
BRAM[39]<= 32'hBF44C130;
BRAM[40]<= 32'h600C6804;
BRAM[41]<= 32'h00004770;
BRAM[42]<= 32'h24002300;
BRAM[43]<= 32'h26002500;
BRAM[44]<= 32'hBF283A10;
BRAM[45]<= 32'hD8FBC178;
BRAM[46]<= 32'hBF280752;
BRAM[47]<= 32'hBF48C130;
BRAM[48]<= 32'h4770600B;
BRAM[49]<= 32'hBD1FB51F;
BRAM[50]<= 32'hBD10B510;
BRAM[51]<= 32'hF892F000;
BRAM[52]<= 32'hF7FF4611;
BRAM[53]<= 32'hF001FFF7;
BRAM[54]<= 32'hF000F9C9;
BRAM[55]<= 32'hB403F8C4;
BRAM[56]<= 32'hFFF2F7FF;
BRAM[57]<= 32'hF001BC03;
BRAM[58]<= 32'h0000F98F;
BRAM[59]<= 32'h4780481E;
BRAM[60]<= 32'h4700481E;
BRAM[61]<= 32'hF001B500;
BRAM[62]<= 32'hBD00F8D5;
BRAM[63]<= 32'hF000B500;
BRAM[64]<= 32'hBD00FA9B;
BRAM[65]<= 32'hF001B500;
BRAM[66]<= 32'hBD00F8CC;
BRAM[67]<= 32'hF000B500;
BRAM[68]<= 32'hBD00F8B7;
BRAM[69]<= 32'hF001B500;
BRAM[70]<= 32'hBD00F976;
BRAM[71]<= 32'hF001B500;
BRAM[72]<= 32'hBD00F906;
BRAM[73]<= 32'hF000B500;
BRAM[74]<= 32'hBD00F8AC;
BRAM[75]<= 32'hF001B500;
BRAM[76]<= 32'hBD00F8FD;
BRAM[77]<= 32'hF001B500;
BRAM[78]<= 32'hBD00F947;
BRAM[79]<= 32'hF001B500;
BRAM[80]<= 32'hBD00F960;
BRAM[81]<= 32'hF001B500;
BRAM[82]<= 32'hBD00F95D;
BRAM[83]<= 32'hF001B500;
BRAM[84]<= 32'hBD00F957;
BRAM[85]<= 32'hF000B500;
BRAM[86]<= 32'hBD00F8A7;
BRAM[87]<= 32'h49054804;
BRAM[88]<= 32'h4B064A05;
BRAM[89]<= 32'h00004770;
BRAM[90]<= 32'h000013CD;
BRAM[91]<= 32'h0000146D;
BRAM[92]<= 32'h20000080;
BRAM[93]<= 32'h2000A080;
BRAM[94]<= 32'h20005080;
BRAM[95]<= 32'h20005080;
BRAM[96]<= 32'h4904B40F;
BRAM[97]<= 32'hAA03B510;
BRAM[98]<= 32'hF0009802;
BRAM[99]<= 32'hBC10F809;
BRAM[100]<= 32'hFB14F85D;
BRAM[101]<= 32'h20000010;
BRAM[102]<= 32'h47704770;
BRAM[103]<= 32'h00004770;
BRAM[104]<= 32'hB5704B07;
BRAM[105]<= 32'h447B460D;
BRAM[106]<= 32'hF811F000;
BRAM[107]<= 32'h46284604;
BRAM[108]<= 32'hF948F001;
BRAM[109]<= 32'hF04FB110;
BRAM[110]<= 32'hBD7030FF;
BRAM[111]<= 32'hBD704620;
BRAM[112]<= 32'h000012A3;
BRAM[113]<= 32'h1C4A6901;
BRAM[114]<= 32'h78086102;
BRAM[115]<= 32'hB5004770;
BRAM[116]<= 32'hE9CDB08F;
BRAM[117]<= 32'h21003101;
BRAM[118]<= 32'h49059105;
BRAM[119]<= 32'hE9CD4479;
BRAM[120]<= 32'h46111003;
BRAM[121]<= 32'hF0004668;
BRAM[122]<= 32'hB00FF82A;
BRAM[123]<= 32'h0000BD00;
BRAM[124]<= 32'hFFFFFFE5;
BRAM[125]<= 32'hF0004675;
BRAM[126]<= 32'h46AEF83F;
BRAM[127]<= 32'h46690005;
BRAM[128]<= 32'hF0204653;
BRAM[129]<= 32'h46850007;
BRAM[130]<= 32'hB520B018;
BRAM[131]<= 32'hFFA6F7FF;
BRAM[132]<= 32'h4020E8BD;
BRAM[133]<= 32'h0600F04F;
BRAM[134]<= 32'h0700F04F;
BRAM[135]<= 32'h0800F04F;
BRAM[136]<= 32'h0B00F04F;
BRAM[137]<= 32'h0107F021;
BRAM[138]<= 32'hE8AC46AC;
BRAM[139]<= 32'hE8AC09C0;
BRAM[140]<= 32'hE8AC09C0;
BRAM[141]<= 32'hE8AC09C0;
BRAM[142]<= 32'h468D09C0;
BRAM[143]<= 32'hE92D4770;
BRAM[144]<= 32'h460641F0;
BRAM[145]<= 32'hE9D62400;
BRAM[146]<= 32'h68F57001;
BRAM[147]<= 32'h46304680;
BRAM[148]<= 32'h4641E003;
BRAM[149]<= 32'h1C6447B8;
BRAM[150]<= 32'h47A84630;
BRAM[151]<= 32'hD1F82800;
BRAM[152]<= 32'hE8BD4620;
BRAM[153]<= 32'hB51081F0;
BRAM[154]<= 32'hF3AF4604;
BRAM[155]<= 32'h46208000;
BRAM[156]<= 32'h4010E8BD;
BRAM[157]<= 32'hBF33F7FF;
BRAM[158]<= 32'h47704800;
BRAM[159]<= 32'h2000001C;
BRAM[160]<= 32'h47704770;
BRAM[161]<= 32'h2003B508;
BRAM[162]<= 32'h0000F88D;
BRAM[163]<= 32'hF88D2002;
BRAM[164]<= 32'h20030001;
BRAM[165]<= 32'h0002F88D;
BRAM[166]<= 32'hF88D2001;
BRAM[167]<= 32'h46680003;
BRAM[168]<= 32'hF802F001;
BRAM[169]<= 32'h0000BD08;
BRAM[170]<= 32'hF44FB510;
BRAM[171]<= 32'hF00170FA;
BRAM[172]<= 32'hF64FF8BF;
BRAM[173]<= 32'hF04F70FF;
BRAM[174]<= 32'h638841A0;
BRAM[175]<= 32'h780048BE;
BRAM[176]<= 32'hD14D2800;
BRAM[177]<= 32'hF0002006;
BRAM[178]<= 32'hB958F998;
BRAM[179]<= 32'h2006BF00;
BRAM[180]<= 32'hF993F000;
BRAM[181]<= 32'hD0FA2800;
BRAM[182]<= 32'h46112200;
BRAM[183]<= 32'hF0002005;
BRAM[184]<= 32'hE164FC7B;
BRAM[185]<= 32'hF0002005;
BRAM[186]<= 32'hB958F988;
BRAM[187]<= 32'h2005BF00;
BRAM[188]<= 32'hF983F000;
BRAM[189]<= 32'hD0FA2800;
BRAM[190]<= 32'h21012200;
BRAM[191]<= 32'hF0002005;
BRAM[192]<= 32'hE154FC6B;
BRAM[193]<= 32'hF0002004;
BRAM[194]<= 32'h2800F978;
BRAM[195]<= 32'hBF00D1E9;
BRAM[196]<= 32'hF0002004;
BRAM[197]<= 32'h2800F972;
BRAM[198]<= 32'h48A8D0FA;
BRAM[199]<= 32'h28017800;
BRAM[200]<= 32'hF000D102;
BRAM[201]<= 32'hE142FDAB;
BRAM[202]<= 32'h780048A4;
BRAM[203]<= 32'hD1022802;
BRAM[204]<= 32'hFDE6F000;
BRAM[205]<= 32'h48A1E13B;
BRAM[206]<= 32'h28037800;
BRAM[207]<= 32'hF000D102;
BRAM[208]<= 32'hE134FE2B;
BRAM[209]<= 32'h7800489D;
BRAM[210]<= 32'hD1022804;
BRAM[211]<= 32'hF828F001;
BRAM[212]<= 32'h489AE12D;
BRAM[213]<= 32'h28057800;
BRAM[214]<= 32'hF001D1C3;
BRAM[215]<= 32'hE126F82B;
BRAM[216]<= 32'h78004895;
BRAM[217]<= 32'hD1372801;
BRAM[218]<= 32'hF0002006;
BRAM[219]<= 32'hB958F946;
BRAM[220]<= 32'h2006BF00;
BRAM[221]<= 32'hF941F000;
BRAM[222]<= 32'hD0FA2800;
BRAM[223]<= 32'h46112200;
BRAM[224]<= 32'hF0002004;
BRAM[225]<= 32'hE112FC29;
BRAM[226]<= 32'hF0002005;
BRAM[227]<= 32'hB958F936;
BRAM[228]<= 32'h2005BF00;
BRAM[229]<= 32'hF931F000;
BRAM[230]<= 32'hD0FA2800;
BRAM[231]<= 32'h21012200;
BRAM[232]<= 32'hF0002004;
BRAM[233]<= 32'hE102FC19;
BRAM[234]<= 32'hF0002004;
BRAM[235]<= 32'h2800F926;
BRAM[236]<= 32'hBF00D197;
BRAM[237]<= 32'hF0002004;
BRAM[238]<= 32'h2800F920;
BRAM[239]<= 32'h487FD0FA;
BRAM[240]<= 32'h28047800;
BRAM[241]<= 32'hF000D102;
BRAM[242]<= 32'hE0F0FC51;
BRAM[243]<= 32'h7800487B;
BRAM[244]<= 32'h497B1E40;
BRAM[245]<= 32'hE0EA7008;
BRAM[246]<= 32'h78004877;
BRAM[247]<= 32'hD1692802;
BRAM[248]<= 32'hF0002006;
BRAM[249]<= 32'hB958F90A;
BRAM[250]<= 32'h2006BF00;
BRAM[251]<= 32'hF905F000;
BRAM[252]<= 32'hD0FA2800;
BRAM[253]<= 32'h46112200;
BRAM[254]<= 32'hF0002005;
BRAM[255]<= 32'hE0D6FBED;
BRAM[256]<= 32'hF0002005;
BRAM[257]<= 32'hB958F8FA;
BRAM[258]<= 32'h2005BF00;
BRAM[259]<= 32'hF8F5F000;
BRAM[260]<= 32'hD0FA2800;
BRAM[261]<= 32'h21012200;
BRAM[262]<= 32'hF0002005;
BRAM[263]<= 32'hE0C6FBDD;
BRAM[264]<= 32'hF0002004;
BRAM[265]<= 32'hB960F8EA;
BRAM[266]<= 32'h2004BF00;
BRAM[267]<= 32'hF8E5F000;
BRAM[268]<= 32'hD0FA2800;
BRAM[269]<= 32'h78004861;
BRAM[270]<= 32'hD1892805;
BRAM[271]<= 32'hFC16F000;
BRAM[272]<= 32'h2003E0B5;
BRAM[273]<= 32'hF8D9F000;
BRAM[274]<= 32'hBF00BB98;
BRAM[275]<= 32'hF0002003;
BRAM[276]<= 32'h2800F8D4;
BRAM[277]<= 32'h4859D0FA;
BRAM[278]<= 32'h28017800;
BRAM[279]<= 32'h4859D10A;
BRAM[280]<= 32'h0A006900;
BRAM[281]<= 32'h49571C40;
BRAM[282]<= 32'hF3606909;
BRAM[283]<= 32'h4855210F;
BRAM[284]<= 32'hE0296101;
BRAM[285]<= 32'h78004851;
BRAM[286]<= 32'hD10A2802;
BRAM[287]<= 32'h69004851;
BRAM[288]<= 32'h1C400C00;
BRAM[289]<= 32'h6909494F;
BRAM[290]<= 32'h4117F360;
BRAM[291]<= 32'h6101484D;
BRAM[292]<= 32'h484AE01A;
BRAM[293]<= 32'h28037800;
BRAM[294]<= 32'h484AD10D;
BRAM[295]<= 32'h21016900;
BRAM[296]<= 32'h6110EB01;
BRAM[297]<= 32'h69004847;
BRAM[298]<= 32'h601FF361;
BRAM[299]<= 32'h61084945;
BRAM[300]<= 32'hE00CE00A;
BRAM[301]<= 32'h4841E050;
BRAM[302]<= 32'h28047800;
BRAM[303]<= 32'h4841D104;
BRAM[304]<= 32'h1C406940;
BRAM[305]<= 32'h6148493F;
BRAM[306]<= 32'hFC2AF000;
BRAM[307]<= 32'h2002E06F;
BRAM[308]<= 32'hF893F000;
BRAM[309]<= 32'hD16A2800;
BRAM[310]<= 32'h2002BF00;
BRAM[311]<= 32'hF88DF000;
BRAM[312]<= 32'hD0FA2800;
BRAM[313]<= 32'h78004835;
BRAM[314]<= 32'hD10A2801;
BRAM[315]<= 32'h69004835;
BRAM[316]<= 32'h1E400A00;
BRAM[317]<= 32'h69094933;
BRAM[318]<= 32'h210FF360;
BRAM[319]<= 32'h61014831;
BRAM[320]<= 32'h482EE027;
BRAM[321]<= 32'h28027800;
BRAM[322]<= 32'h482ED10A;
BRAM[323]<= 32'h0C006900;
BRAM[324]<= 32'h492C1E40;
BRAM[325]<= 32'hF3606909;
BRAM[326]<= 32'h482A4117;
BRAM[327]<= 32'hE0186101;
BRAM[328]<= 32'h78004826;
BRAM[329]<= 32'hD10B2803;
BRAM[330]<= 32'h69004826;
BRAM[331]<= 32'hEBC12101;
BRAM[332]<= 32'h48246110;
BRAM[333]<= 32'hF3616900;
BRAM[334]<= 32'h4922601F;
BRAM[335]<= 32'hE0086108;
BRAM[336]<= 32'h7800481E;
BRAM[337]<= 32'hD1042804;
BRAM[338]<= 32'h6940481E;
BRAM[339]<= 32'h491D1E40;
BRAM[340]<= 32'hF0006148;
BRAM[341]<= 32'hE02AFBE5;
BRAM[342]<= 32'h78004817;
BRAM[343]<= 32'hD1262803;
BRAM[344]<= 32'hF0002004;
BRAM[345]<= 32'hB948F84A;
BRAM[346]<= 32'h2004BF00;
BRAM[347]<= 32'hF845F000;
BRAM[348]<= 32'hD0FA2800;
BRAM[349]<= 32'h49142001;
BRAM[350]<= 32'hE0187008;
BRAM[351]<= 32'hF0002003;
BRAM[352]<= 32'hB940F83C;
BRAM[353]<= 32'h2003BF00;
BRAM[354]<= 32'hF837F000;
BRAM[355]<= 32'hD0FA2800;
BRAM[356]<= 32'hFF06F000;
BRAM[357]<= 32'h2002E00B;
BRAM[358]<= 32'hF82FF000;
BRAM[359]<= 32'hBF00B938;
BRAM[360]<= 32'hF0002002;
BRAM[361]<= 32'h2800F82A;
BRAM[362]<= 32'hF000D0FA;
BRAM[363]<= 32'hA007FF03;
BRAM[364]<= 32'hFDE6F7FF;
BRAM[365]<= 32'h0000BD10;
BRAM[366]<= 32'h2000000D;
BRAM[367]<= 32'h2000000E;
BRAM[368]<= 32'h2000000C;
BRAM[369]<= 32'h40001000;
BRAM[370]<= 32'h2000000F;
BRAM[371]<= 32'h4F495047;
BRAM[372]<= 32'h00000A21;
BRAM[373]<= 32'h7083F64F;
BRAM[374]<= 32'h41A0F04F;
BRAM[375]<= 32'h207C6108;
BRAM[376]<= 32'h20006148;
BRAM[377]<= 32'hF64F6188;
BRAM[378]<= 32'h61C870FF;
BRAM[379]<= 32'h207C6048;
BRAM[380]<= 32'hF64F6208;
BRAM[381]<= 32'h634870FF;
BRAM[382]<= 32'h46014770;
BRAM[383]<= 32'h40A0F04F;
BRAM[384]<= 32'h40C86800;
BRAM[385]<= 32'h0001F000;
BRAM[386]<= 32'hB9494770;
BRAM[387]<= 32'h42A0F04F;
BRAM[388]<= 32'h23016852;
BRAM[389]<= 32'h439A4083;
BRAM[390]<= 32'h43A0F04F;
BRAM[391]<= 32'hE00A605A;
BRAM[392]<= 32'hD1082901;
BRAM[393]<= 32'h42A0F04F;
BRAM[394]<= 32'h23016852;
BRAM[395]<= 32'h431A4083;
BRAM[396]<= 32'h43A0F04F;
BRAM[397]<= 32'h4770605A;
BRAM[398]<= 32'hA002B510;
BRAM[399]<= 32'hFDA0F7FF;
BRAM[400]<= 32'h0000BD10;
BRAM[401]<= 32'h64726148;
BRAM[402]<= 32'h6C756146;
BRAM[403]<= 32'h000A2174;
BRAM[404]<= 32'h41F0E92D;
BRAM[405]<= 32'h460D4604;
BRAM[406]<= 32'h461F4616;
BRAM[407]<= 32'hF000202A;
BRAM[408]<= 32'hF3C4FA6F;
BRAM[409]<= 32'hF0002007;
BRAM[410]<= 32'hB2E0FA61;
BRAM[411]<= 32'hFA5EF000;
BRAM[412]<= 32'h2007F3C6;
BRAM[413]<= 32'hFA5AF000;
BRAM[414]<= 32'hF000B2F0;
BRAM[415]<= 32'h202BFA57;
BRAM[416]<= 32'hFA5EF000;
BRAM[417]<= 32'h2007F3C5;
BRAM[418]<= 32'hFA50F000;
BRAM[419]<= 32'hF000B2E8;
BRAM[420]<= 32'hF3C7FA4D;
BRAM[421]<= 32'hF0002007;
BRAM[422]<= 32'hB2F8FA49;
BRAM[423]<= 32'hFA46F000;
BRAM[424]<= 32'hF000202C;
BRAM[425]<= 32'hE8BDFA4D;
BRAM[426]<= 32'hB57081F0;
BRAM[427]<= 32'hF2404606;
BRAM[428]<= 32'hF240133F;
BRAM[429]<= 32'h210012DF;
BRAM[430]<= 32'hF7FF4608;
BRAM[431]<= 32'h2400FFC9;
BRAM[432]<= 32'h2500E009;
BRAM[433]<= 32'h4630E003;
BRAM[434]<= 32'hFA1EF000;
BRAM[435]<= 32'hF5B51C6D;
BRAM[436]<= 32'hD3F87FA0;
BRAM[437]<= 32'hF5B41C64;
BRAM[438]<= 32'hD3F27FF0;
BRAM[439]<= 32'hE92DBD70;
BRAM[440]<= 32'hB0854FFF;
BRAM[441]<= 32'h468A4681;
BRAM[442]<= 32'h90032000;
BRAM[443]<= 32'h98074683;
BRAM[444]<= 32'h0409EBA0;
BRAM[445]<= 32'hEBA09808;
BRAM[446]<= 32'hF8CD060A;
BRAM[447]<= 32'hF8CD9008;
BRAM[448]<= 32'h2C00A004;
BRAM[449]<= 32'h2701DD01;
BRAM[450]<= 32'hB90CE005;
BRAM[451]<= 32'hE0022700;
BRAM[452]<= 32'h37FFF04F;
BRAM[453]<= 32'h2E004264;
BRAM[454]<= 32'hF04FDD02;
BRAM[455]<= 32'hE0060801;
BRAM[456]<= 32'hF04FB916;
BRAM[457]<= 32'hE0020800;
BRAM[458]<= 32'h38FFF04F;
BRAM[459]<= 32'h42B44266;
BRAM[460]<= 32'h4625DD01;
BRAM[461]<= 32'h4635E000;
BRAM[462]<= 32'h90042000;
BRAM[463]<= 32'h9A12E01B;
BRAM[464]<= 32'h1001E9DD;
BRAM[465]<= 32'hF81EF000;
BRAM[466]<= 32'h44209803;
BRAM[467]<= 32'h44B39003;
BRAM[468]<= 32'h42A89803;
BRAM[469]<= 32'h9803DD05;
BRAM[470]<= 32'h90031B40;
BRAM[471]<= 32'h44389802;
BRAM[472]<= 32'h45AB9002;
BRAM[473]<= 32'hEBABDD04;
BRAM[474]<= 32'h98010B05;
BRAM[475]<= 32'h90014440;
BRAM[476]<= 32'h1C409804;
BRAM[477]<= 32'h1C699004;
BRAM[478]<= 32'h42889804;
BRAM[479]<= 32'hB009D3DF;
BRAM[480]<= 32'h8FF0E8BD;
BRAM[481]<= 32'h4604B570;
BRAM[482]<= 32'h4616460D;
BRAM[483]<= 32'h4622462B;
BRAM[484]<= 32'h46204629;
BRAM[485]<= 32'hFF5CF7FF;
BRAM[486]<= 32'hF0004630;
BRAM[487]<= 32'hBD70F9B5;
BRAM[488]<= 32'h43F8E92D;
BRAM[489]<= 32'h460E4605;
BRAM[490]<= 32'h46984617;
BRAM[491]<= 32'h46339C08;
BRAM[492]<= 32'h4631463A;
BRAM[493]<= 32'h94004628;
BRAM[494]<= 32'hFF91F7FF;
BRAM[495]<= 32'h462A4643;
BRAM[496]<= 32'h46284631;
BRAM[497]<= 32'hF7FF9400;
BRAM[498]<= 32'h4643FF8A;
BRAM[499]<= 32'h4641463A;
BRAM[500]<= 32'h94004628;
BRAM[501]<= 32'hFF83F7FF;
BRAM[502]<= 32'h463A4643;
BRAM[503]<= 32'h46384631;
BRAM[504]<= 32'hF7FF9400;
BRAM[505]<= 32'hE8BDFF7C;
BRAM[506]<= 32'h000083F8;
BRAM[507]<= 32'h5FF0E92D;
BRAM[508]<= 32'h46894605;
BRAM[509]<= 32'h461E4693;
BRAM[510]<= 32'hA028F8DD;
BRAM[511]<= 32'hE0322400;
BRAM[512]<= 32'h0106EB09;
BRAM[513]<= 32'hEB041E4B;
BRAM[514]<= 32'hEB050144;
BRAM[515]<= 32'h443101C1;
BRAM[516]<= 32'hEB041E4A;
BRAM[517]<= 32'hEB050144;
BRAM[518]<= 32'h464900C1;
BRAM[519]<= 32'hFF18F7FF;
BRAM[520]<= 32'h0800F04F;
BRAM[521]<= 32'h2700E01A;
BRAM[522]<= 32'hEB04E012;
BRAM[523]<= 32'hEB0800C4;
BRAM[524]<= 32'h490F00C0;
BRAM[525]<= 32'h21015C08;
BRAM[526]<= 32'h400840B9;
BRAM[527]<= 32'h4650B118;
BRAM[528]<= 32'hF962F000;
BRAM[529]<= 32'h480BE002;
BRAM[530]<= 32'hF95EF000;
BRAM[531]<= 32'hB2C71C78;
BRAM[532]<= 32'hDBEA2F08;
BRAM[533]<= 32'h0001F108;
BRAM[534]<= 32'h08FFF000;
BRAM[535]<= 32'h0F48F1B8;
BRAM[536]<= 32'h1C60DBE1;
BRAM[537]<= 32'h2C07B2C4;
BRAM[538]<= 32'hE8BDDBCA;
BRAM[539]<= 32'h00009FF0;
BRAM[540]<= 32'h00001C04;
BRAM[541]<= 32'h00FCFCFC;
BRAM[542]<= 32'h5FF0E92D;
BRAM[543]<= 32'h468B4607;
BRAM[544]<= 32'h469A4691;
BRAM[545]<= 32'h09C7F107;
BRAM[546]<= 32'h0A95F10B;
BRAM[547]<= 32'h464A4653;
BRAM[548]<= 32'h46384659;
BRAM[549]<= 32'hFEDCF7FF;
BRAM[550]<= 32'hE03B2400;
BRAM[551]<= 32'hF8104855;
BRAM[552]<= 32'h25038004;
BRAM[553]<= 32'h0068E033;
BRAM[554]<= 32'hF000FA48;
BRAM[555]<= 32'h0603F000;
BRAM[556]<= 32'h20FFB94E;
BRAM[557]<= 32'hF93AF000;
BRAM[558]<= 32'hF0002000;
BRAM[559]<= 32'h2000F937;
BRAM[560]<= 32'hF934F000;
BRAM[561]<= 32'h2E01E022;
BRAM[562]<= 32'h20FFD109;
BRAM[563]<= 32'hF92EF000;
BRAM[564]<= 32'hF0002000;
BRAM[565]<= 32'h2000F92B;
BRAM[566]<= 32'hF928F000;
BRAM[567]<= 32'h2E02E016;
BRAM[568]<= 32'h2000D109;
BRAM[569]<= 32'hF922F000;
BRAM[570]<= 32'hF000205C;
BRAM[571]<= 32'h20E4F91F;
BRAM[572]<= 32'hF91CF000;
BRAM[573]<= 32'h2E03E00A;
BRAM[574]<= 32'h20FFD108;
BRAM[575]<= 32'hF916F000;
BRAM[576]<= 32'hF00020FF;
BRAM[577]<= 32'h20FFF913;
BRAM[578]<= 32'hF910F000;
BRAM[579]<= 32'h2D001E6D;
BRAM[580]<= 32'h1C64DAC9;
BRAM[581]<= 32'h504CF641;
BRAM[582]<= 32'hDBBF4284;
BRAM[583]<= 32'h0109EB07;
BRAM[584]<= 32'hEBC32378;
BRAM[585]<= 32'hF1010151;
BRAM[586]<= 32'hEB0702EF;
BRAM[587]<= 32'hEBC30109;
BRAM[588]<= 32'hF10A0051;
BRAM[589]<= 32'hF10A0322;
BRAM[590]<= 32'hF7FF010A;
BRAM[591]<= 32'h2400FE89;
BRAM[592]<= 32'h482DE022;
BRAM[593]<= 32'h8004F810;
BRAM[594]<= 32'hE01A2507;
BRAM[595]<= 32'hF005FA48;
BRAM[596]<= 32'h0601F000;
BRAM[597]<= 32'h20FFB94E;
BRAM[598]<= 32'hF8E8F000;
BRAM[599]<= 32'hF00020FF;
BRAM[600]<= 32'h20FFF8E5;
BRAM[601]<= 32'hF8E2F000;
BRAM[602]<= 32'h2E01E00A;
BRAM[603]<= 32'h2000D108;
BRAM[604]<= 32'hF8DCF000;
BRAM[605]<= 32'hF0002000;
BRAM[606]<= 32'h2000F8D9;
BRAM[607]<= 32'hF8D6F000;
BRAM[608]<= 32'h2D001E6D;
BRAM[609]<= 32'h1C64DAE2;
BRAM[610]<= 32'h20EEF240;
BRAM[611]<= 32'hDBD84284;
BRAM[612]<= 32'hF2402329;
BRAM[613]<= 32'h210A128F;
BRAM[614]<= 32'hF7FF2050;
BRAM[615]<= 32'h2400FE59;
BRAM[616]<= 32'h4816E022;
BRAM[617]<= 32'h8004F810;
BRAM[618]<= 32'hE01A2507;
BRAM[619]<= 32'hF005FA48;
BRAM[620]<= 32'h0601F000;
BRAM[621]<= 32'h20FFB94E;
BRAM[622]<= 32'hF8B8F000;
BRAM[623]<= 32'hF00020FF;
BRAM[624]<= 32'h20FFF8B5;
BRAM[625]<= 32'hF8B2F000;
BRAM[626]<= 32'h2E01E00A;
BRAM[627]<= 32'h20FFD108;
BRAM[628]<= 32'hF8ACF000;
BRAM[629]<= 32'hF0002000;
BRAM[630]<= 32'h2000F8A9;
BRAM[631]<= 32'hF8A6F000;
BRAM[632]<= 32'h2D001E6D;
BRAM[633]<= 32'h1C64DAE2;
BRAM[634]<= 32'h6FA0F5B4;
BRAM[635]<= 32'hE8BDDBD9;
BRAM[636]<= 32'h00009FF0;
BRAM[637]<= 32'h0000273C;
BRAM[638]<= 32'h00004488;
BRAM[639]<= 32'h0000223C;
BRAM[640]<= 32'h5FF0E92D;
BRAM[641]<= 32'h46894606;
BRAM[642]<= 32'h469A4615;
BRAM[643]<= 32'hE0722400;
BRAM[644]<= 32'h030FF109;
BRAM[645]<= 32'h01C4EB06;
BRAM[646]<= 32'hEB061DCA;
BRAM[647]<= 32'h464900C4;
BRAM[648]<= 32'hFE16F7FF;
BRAM[649]<= 32'h28305D28;
BRAM[650]<= 32'h5D28DB08;
BRAM[651]<= 32'hDC052839;
BRAM[652]<= 32'h38305D28;
BRAM[653]<= 32'hEB012100;
BRAM[654]<= 32'hE03B1B00;
BRAM[655]<= 32'h28415D28;
BRAM[656]<= 32'h5D28DB08;
BRAM[657]<= 32'hDC05285A;
BRAM[658]<= 32'h38415D28;
BRAM[659]<= 32'hEB0121A0;
BRAM[660]<= 32'hE02F1B00;
BRAM[661]<= 32'h28615D28;
BRAM[662]<= 32'h5D28DB09;
BRAM[663]<= 32'hDC06287A;
BRAM[664]<= 32'h38615D28;
BRAM[665]<= 32'h7110F44F;
BRAM[666]<= 32'h1B00EB01;
BRAM[667]<= 32'h5D28E022;
BRAM[668]<= 32'hD102285F;
BRAM[669]<= 32'h7B78F44F;
BRAM[670]<= 32'h5D28E01C;
BRAM[671]<= 32'hD102283A;
BRAM[672]<= 32'h7B7CF44F;
BRAM[673]<= 32'h5D28E016;
BRAM[674]<= 32'hD102283C;
BRAM[675]<= 32'h6B80F44F;
BRAM[676]<= 32'h5D28E010;
BRAM[677]<= 32'hD1022820;
BRAM[678]<= 32'h6B82F44F;
BRAM[679]<= 32'h5D28E00A;
BRAM[680]<= 32'hD102282B;
BRAM[681]<= 32'h6B84F44F;
BRAM[682]<= 32'h5D28E004;
BRAM[683]<= 32'hD101282D;
BRAM[684]<= 32'h6B86F44F;
BRAM[685]<= 32'h0800F04F;
BRAM[686]<= 32'h2700E018;
BRAM[687]<= 32'hEB0BE010;
BRAM[688]<= 32'h490F0008;
BRAM[689]<= 32'h21015C08;
BRAM[690]<= 32'h400840B9;
BRAM[691]<= 32'h4650B118;
BRAM[692]<= 32'hF81AF000;
BRAM[693]<= 32'h480BE002;
BRAM[694]<= 32'hF816F000;
BRAM[695]<= 32'hB2C71C78;
BRAM[696]<= 32'hDBEC2F08;
BRAM[697]<= 32'h0001F108;
BRAM[698]<= 32'h08FFF000;
BRAM[699]<= 32'h0F10F1B8;
BRAM[700]<= 32'h1C60DBE3;
BRAM[701]<= 32'h5D28B2C4;
BRAM[702]<= 32'hD1892800;
BRAM[703]<= 32'h9FF0E8BD;
BRAM[704]<= 32'h00001DFC;
BRAM[705]<= 32'h00FCFCFC;
BRAM[706]<= 32'h4604B510;
BRAM[707]<= 32'h200F2101;
BRAM[708]<= 32'hFD7BF7FF;
BRAM[709]<= 32'h4007F3C4;
BRAM[710]<= 32'hF81CF000;
BRAM[711]<= 32'h2007F3C4;
BRAM[712]<= 32'hF818F000;
BRAM[713]<= 32'hF000B2E0;
BRAM[714]<= 32'hBD10F815;
BRAM[715]<= 32'h4604B510;
BRAM[716]<= 32'h200F2101;
BRAM[717]<= 32'hFD69F7FF;
BRAM[718]<= 32'hF0004620;
BRAM[719]<= 32'hBD10F80B;
BRAM[720]<= 32'h4604B510;
BRAM[721]<= 32'h200F2100;
BRAM[722]<= 32'hFD5FF7FF;
BRAM[723]<= 32'hF0004620;
BRAM[724]<= 32'hBD10F801;
BRAM[725]<= 32'h4604B570;
BRAM[726]<= 32'hE0172500;
BRAM[727]<= 32'h200C2100;
BRAM[728]<= 32'hFD53F7FF;
BRAM[729]<= 32'h0080F004;
BRAM[730]<= 32'h2101B120;
BRAM[731]<= 32'hF7FF200D;
BRAM[732]<= 32'hE003FD4C;
BRAM[733]<= 32'h200D2100;
BRAM[734]<= 32'hFD47F7FF;
BRAM[735]<= 32'h200C2101;
BRAM[736]<= 32'hFD43F7FF;
BRAM[737]<= 32'h0E040660;
BRAM[738]<= 32'hB2C51C68;
BRAM[739]<= 32'hDBE52D08;
BRAM[740]<= 32'h0000BD70;
BRAM[741]<= 32'h2400B510;
BRAM[742]<= 32'hEB04E00C;
BRAM[743]<= 32'h00C00044;
BRAM[744]<= 32'h0178F100;
BRAM[745]<= 32'hA2064B05;
BRAM[746]<= 32'h7091F44F;
BRAM[747]<= 32'hFF28F7FF;
BRAM[748]<= 32'hB2C41C60;
BRAM[749]<= 32'hDBF02C0A;
BRAM[750]<= 32'h0000BD10;
BRAM[751]<= 32'h00FCFCFC;
BRAM[752]<= 32'h20202020;
BRAM[753]<= 32'h20202020;
BRAM[754]<= 32'h20202020;
BRAM[755]<= 32'h20202020;
BRAM[756]<= 32'h20202020;
BRAM[757]<= 32'h00002020;
BRAM[758]<= 32'h4604B570;
BRAM[759]<= 32'h4616460D;
BRAM[760]<= 32'h7800481F;
BRAM[761]<= 32'hEB001E40;
BRAM[762]<= 32'h00C00040;
BRAM[763]<= 32'h0178F100;
BRAM[764]<= 32'hA21C2300;
BRAM[765]<= 32'h70D9F44F;
BRAM[766]<= 32'hFF02F7FF;
BRAM[767]<= 32'h2D01BB46;
BRAM[768]<= 32'h4817D105;
BRAM[769]<= 32'h1C407800;
BRAM[770]<= 32'h70084915;
BRAM[771]<= 32'h4814E004;
BRAM[772]<= 32'h1E407800;
BRAM[773]<= 32'h70084912;
BRAM[774]<= 32'h78004811;
BRAM[775]<= 32'hDD0242A0;
BRAM[776]<= 32'h490F2001;
BRAM[777]<= 32'h480E7008;
BRAM[778]<= 32'h28007800;
BRAM[779]<= 32'h480CDC01;
BRAM[780]<= 32'h480B7004;
BRAM[781]<= 32'h1E407800;
BRAM[782]<= 32'h0040EB00;
BRAM[783]<= 32'hF10000C0;
BRAM[784]<= 32'h23000178;
BRAM[785]<= 32'hF44FA208;
BRAM[786]<= 32'hF7FF70D9;
BRAM[787]<= 32'hE006FED9;
BRAM[788]<= 32'hA2052300;
BRAM[789]<= 32'hF44F2178;
BRAM[790]<= 32'hF7FF70D9;
BRAM[791]<= 32'hBD70FED1;
BRAM[792]<= 32'h2000000E;
BRAM[793]<= 32'h00000020;
BRAM[794]<= 32'h0000003C;
BRAM[795]<= 32'h2000B510;
BRAM[796]<= 32'h70084917;
BRAM[797]<= 32'hFF8EF7FF;
BRAM[798]<= 32'h21002201;
BRAM[799]<= 32'hF7FF2005;
BRAM[800]<= 32'h2001FFAB;
BRAM[801]<= 32'h70084913;
BRAM[802]<= 32'hA2132300;
BRAM[803]<= 32'hF44F2178;
BRAM[804]<= 32'hF7FF7091;
BRAM[805]<= 32'h2300FEB5;
BRAM[806]<= 32'h2190A212;
BRAM[807]<= 32'h7091F44F;
BRAM[808]<= 32'hFEAEF7FF;
BRAM[809]<= 32'hA2122300;
BRAM[810]<= 32'hF44F21A8;
BRAM[811]<= 32'hF7FF7091;
BRAM[812]<= 32'h2300FEA7;
BRAM[813]<= 32'h21C0A212;
BRAM[814]<= 32'h7091F44F;
BRAM[815]<= 32'hFEA0F7FF;
BRAM[816]<= 32'hA2132300;
BRAM[817]<= 32'hF44F21D8;
BRAM[818]<= 32'hF7FF7091;
BRAM[819]<= 32'hBD10FE99;
BRAM[820]<= 32'h2000000D;
BRAM[821]<= 32'h2000000E;
BRAM[822]<= 32'h2044454C;
BRAM[823]<= 32'h65646F6D;
BRAM[824]<= 32'h00003A6C;
BRAM[825]<= 32'h20737953;
BRAM[826]<= 32'h3A746573;
BRAM[827]<= 32'h00000000;
BRAM[828]<= 32'h20737953;
BRAM[829]<= 32'h696E6F6D;
BRAM[830]<= 32'h3A726F74;
BRAM[831]<= 32'h00000000;
BRAM[832]<= 32'h65636341;
BRAM[833]<= 32'h6172656C;
BRAM[834]<= 32'h20726F74;
BRAM[835]<= 32'h00545352;
BRAM[836]<= 32'h65636341;
BRAM[837]<= 32'h6172656C;
BRAM[838]<= 32'h20726F74;
BRAM[839]<= 32'h004E5552;
BRAM[840]<= 32'h2001B51C;
BRAM[841]<= 32'hFB04F000;
BRAM[842]<= 32'h20644604;
BRAM[843]<= 32'hF0F0FBB4;
BRAM[844]<= 32'hB2C03030;
BRAM[845]<= 32'h0000F88D;
BRAM[846]<= 32'hFBB42064;
BRAM[847]<= 32'hFB00F1F0;
BRAM[848]<= 32'h210A4011;
BRAM[849]<= 32'hF0F1FBB0;
BRAM[850]<= 32'hF88D3030;
BRAM[851]<= 32'h20640001;
BRAM[852]<= 32'hF1F0FBB4;
BRAM[853]<= 32'h4011FB00;
BRAM[854]<= 32'hFBB0210A;
BRAM[855]<= 32'hFB01F2F1;
BRAM[856]<= 32'h30300012;
BRAM[857]<= 32'h0002F88D;
BRAM[858]<= 32'hF88D2000;
BRAM[859]<= 32'h23000003;
BRAM[860]<= 32'h2178466A;
BRAM[861]<= 32'h70C1F44F;
BRAM[862]<= 32'hFE42F7FF;
BRAM[863]<= 32'hF0002002;
BRAM[864]<= 32'h4604FAD7;
BRAM[865]<= 32'hFBB42064;
BRAM[866]<= 32'h3030F0F0;
BRAM[867]<= 32'hF88DB2C0;
BRAM[868]<= 32'h20640000;
BRAM[869]<= 32'hF1F0FBB4;
BRAM[870]<= 32'h4011FB00;
BRAM[871]<= 32'hFBB0210A;
BRAM[872]<= 32'h3030F0F1;
BRAM[873]<= 32'h0001F88D;
BRAM[874]<= 32'hFBB42064;
BRAM[875]<= 32'hFB00F1F0;
BRAM[876]<= 32'h210A4011;
BRAM[877]<= 32'hF2F1FBB0;
BRAM[878]<= 32'h0012FB01;
BRAM[879]<= 32'hF88D3030;
BRAM[880]<= 32'h23000002;
BRAM[881]<= 32'h2190466A;
BRAM[882]<= 32'h70C1F44F;
BRAM[883]<= 32'hFE18F7FF;
BRAM[884]<= 32'hF0002003;
BRAM[885]<= 32'h4604FAAD;
BRAM[886]<= 32'hFBB42064;
BRAM[887]<= 32'h3030F0F0;
BRAM[888]<= 32'hF88DB2C0;
BRAM[889]<= 32'h20640000;
BRAM[890]<= 32'hF1F0FBB4;
BRAM[891]<= 32'h4011FB00;
BRAM[892]<= 32'hFBB0210A;
BRAM[893]<= 32'h3030F0F1;
BRAM[894]<= 32'h0001F88D;
BRAM[895]<= 32'hFBB42064;
BRAM[896]<= 32'hFB00F1F0;
BRAM[897]<= 32'h210A4011;
BRAM[898]<= 32'hF2F1FBB0;
BRAM[899]<= 32'h0012FB01;
BRAM[900]<= 32'hF88D3030;
BRAM[901]<= 32'h23000002;
BRAM[902]<= 32'h21A8466A;
BRAM[903]<= 32'h70C1F44F;
BRAM[904]<= 32'hFDEEF7FF;
BRAM[905]<= 32'hF0002004;
BRAM[906]<= 32'h4604FA83;
BRAM[907]<= 32'hFBB42064;
BRAM[908]<= 32'h3030F0F0;
BRAM[909]<= 32'hF88DB2C0;
BRAM[910]<= 32'h20640000;
BRAM[911]<= 32'hF1F0FBB4;
BRAM[912]<= 32'h4011FB00;
BRAM[913]<= 32'hFBB0210A;
BRAM[914]<= 32'h3030F0F1;
BRAM[915]<= 32'h0001F88D;
BRAM[916]<= 32'hFBB42064;
BRAM[917]<= 32'hFB00F1F0;
BRAM[918]<= 32'h210A4011;
BRAM[919]<= 32'hF2F1FBB0;
BRAM[920]<= 32'h0012FB01;
BRAM[921]<= 32'hF88D3030;
BRAM[922]<= 32'h23000002;
BRAM[923]<= 32'h21C0466A;
BRAM[924]<= 32'h70C1F44F;
BRAM[925]<= 32'hFDC4F7FF;
BRAM[926]<= 32'h0000BD1C;
BRAM[927]<= 32'h2001B510;
BRAM[928]<= 32'h70084914;
BRAM[929]<= 32'hFE86F7FF;
BRAM[930]<= 32'h21002201;
BRAM[931]<= 32'hF7FF2003;
BRAM[932]<= 32'h2001FEA3;
BRAM[933]<= 32'h70084910;
BRAM[934]<= 32'hA2102300;
BRAM[935]<= 32'hF44F2178;
BRAM[936]<= 32'hF7FF7091;
BRAM[937]<= 32'h2300FDAD;
BRAM[938]<= 32'h2190A20F;
BRAM[939]<= 32'h7091F44F;
BRAM[940]<= 32'hFDA6F7FF;
BRAM[941]<= 32'hA20F2300;
BRAM[942]<= 32'hF44F21A8;
BRAM[943]<= 32'hF7FF7091;
BRAM[944]<= 32'h2300FD9F;
BRAM[945]<= 32'h21C0A20C;
BRAM[946]<= 32'h7091F44F;
BRAM[947]<= 32'hFD98F7FF;
BRAM[948]<= 32'h0000BD10;
BRAM[949]<= 32'h2000000D;
BRAM[950]<= 32'h2000000E;
BRAM[951]<= 32'h7466654C;
BRAM[952]<= 32'h6C6F7220;
BRAM[953]<= 32'h0000006C;
BRAM[954]<= 32'h68676952;
BRAM[955]<= 32'h6F722074;
BRAM[956]<= 32'h00006C6C;
BRAM[957]<= 32'h006C6C41;
BRAM[958]<= 32'h6B636142;
BRAM[959]<= 32'h00000000;
BRAM[960]<= 32'h2002B510;
BRAM[961]<= 32'h70084918;
BRAM[962]<= 32'hFE44F7FF;
BRAM[963]<= 32'h21002201;
BRAM[964]<= 32'hF7FF2005;
BRAM[965]<= 32'h2001FE61;
BRAM[966]<= 32'h70084914;
BRAM[967]<= 32'hA2142300;
BRAM[968]<= 32'hF44F2178;
BRAM[969]<= 32'hF7FF7091;
BRAM[970]<= 32'h2300FD6B;
BRAM[971]<= 32'h2190A211;
BRAM[972]<= 32'h7091F44F;
BRAM[973]<= 32'hFD64F7FF;
BRAM[974]<= 32'hA20F2300;
BRAM[975]<= 32'hF44F21A8;
BRAM[976]<= 32'hF7FF7091;
BRAM[977]<= 32'h2300FD5D;
BRAM[978]<= 32'h21C0A20E;
BRAM[979]<= 32'h7091F44F;
BRAM[980]<= 32'hFD56F7FF;
BRAM[981]<= 32'hA20E2300;
BRAM[982]<= 32'hF44F21D8;
BRAM[983]<= 32'hF7FF7091;
BRAM[984]<= 32'hF7FFFD4F;
BRAM[985]<= 32'hBD10FEDD;
BRAM[986]<= 32'h2000000D;
BRAM[987]<= 32'h2000000E;
BRAM[988]<= 32'h003A2B59;
BRAM[989]<= 32'h003A2D59;
BRAM[990]<= 32'h65726854;
BRAM[991]<= 32'h6C6F6873;
BRAM[992]<= 32'h00003A64;
BRAM[993]<= 32'h70656542;
BRAM[994]<= 32'h6D697420;
BRAM[995]<= 32'h00003A65;
BRAM[996]<= 32'h6B636142;
BRAM[997]<= 32'h00000000;
BRAM[998]<= 32'h2003B510;
BRAM[999]<= 32'h70084920;
BRAM[1000]<= 32'h49202001;
BRAM[1001]<= 32'hF7FF7008;
BRAM[1002]<= 32'h2300FDF5;
BRAM[1003]<= 32'h2178A21E;
BRAM[1004]<= 32'h7091F44F;
BRAM[1005]<= 32'hFD24F7FF;
BRAM[1006]<= 32'hA21E2300;
BRAM[1007]<= 32'hF44F2190;
BRAM[1008]<= 32'hF7FF7091;
BRAM[1009]<= 32'h2300FD1D;
BRAM[1010]<= 32'h21A8A220;
BRAM[1011]<= 32'h7091F44F;
BRAM[1012]<= 32'hFD16F7FF;
BRAM[1013]<= 32'hA2232300;
BRAM[1014]<= 32'hF44F21C0;
BRAM[1015]<= 32'hF7FF7091;
BRAM[1016]<= 32'h2300FD0F;
BRAM[1017]<= 32'h21D8A225;
BRAM[1018]<= 32'h7091F44F;
BRAM[1019]<= 32'hFD08F7FF;
BRAM[1020]<= 32'hA2282300;
BRAM[1021]<= 32'hF44F21F0;
BRAM[1022]<= 32'hF7FF7091;
BRAM[1023]<= 32'h2300FD01;
BRAM[1024]<= 32'hF44FA22A;
BRAM[1025]<= 32'hF44F7184;
BRAM[1026]<= 32'hF7FF7091;
BRAM[1027]<= 32'h2300FCF9;
BRAM[1028]<= 32'hF44FA22C;
BRAM[1029]<= 32'h1C887190;
BRAM[1030]<= 32'hFCF2F7FF;
BRAM[1031]<= 32'h0000BD10;
BRAM[1032]<= 32'h2000000D;
BRAM[1033]<= 32'h2000000E;
BRAM[1034]<= 32'h6F6C6341;
BRAM[1035]<= 32'h74532072;
BRAM[1036]<= 32'h00003A61;
BRAM[1037]<= 32'h20687445;
BRAM[1038]<= 32'h65657073;
BRAM[1039]<= 32'h20203A64;
BRAM[1040]<= 32'h20202020;
BRAM[1041]<= 32'h624B2020;
BRAM[1042]<= 32'h00007370;
BRAM[1043]<= 32'h646C6156;
BRAM[1044]<= 32'h70732061;
BRAM[1045]<= 32'h3A646565;
BRAM[1046]<= 32'h20202020;
BRAM[1047]<= 32'h624B2020;
BRAM[1048]<= 32'h00007370;
BRAM[1049]<= 32'h6D617246;
BRAM[1050]<= 32'h70732065;
BRAM[1051]<= 32'h3A646565;
BRAM[1052]<= 32'h20202020;
BRAM[1053]<= 32'h70662020;
BRAM[1054]<= 32'h00000073;
BRAM[1055]<= 32'h726F7453;
BRAM[1056]<= 32'h70732065;
BRAM[1057]<= 32'h3A646565;
BRAM[1058]<= 32'h20202020;
BRAM[1059]<= 32'h70662020;
BRAM[1060]<= 32'h00000073;
BRAM[1061]<= 32'h20687445;
BRAM[1062]<= 32'h73756472;
BRAM[1063]<= 32'h3A776465;
BRAM[1064]<= 32'h20202020;
BRAM[1065]<= 32'h79422020;
BRAM[1066]<= 32'h00006574;
BRAM[1067]<= 32'h20636556;
BRAM[1068]<= 32'h73756472;
BRAM[1069]<= 32'h3A776465;
BRAM[1070]<= 32'h20202020;
BRAM[1071]<= 32'h79422020;
BRAM[1072]<= 32'h00006574;
BRAM[1073]<= 32'h20414756;
BRAM[1074]<= 32'h73756472;
BRAM[1075]<= 32'h3A776465;
BRAM[1076]<= 32'h20202020;
BRAM[1077]<= 32'h79422020;
BRAM[1078]<= 32'h00006574;
BRAM[1079]<= 32'h2100B510;
BRAM[1080]<= 32'hF7FF200E;
BRAM[1081]<= 32'h20C8FA92;
BRAM[1082]<= 32'hF9A2F000;
BRAM[1083]<= 32'h200E2101;
BRAM[1084]<= 32'hFA8BF7FF;
BRAM[1085]<= 32'hF0002014;
BRAM[1086]<= 32'h2101F99B;
BRAM[1087]<= 32'hF7FF2000;
BRAM[1088]<= 32'h2011FA84;
BRAM[1089]<= 32'hFD1CF7FF;
BRAM[1090]<= 32'hF000203C;
BRAM[1091]<= 32'h20F2F991;
BRAM[1092]<= 32'hFD16F7FF;
BRAM[1093]<= 32'hF7FF2018;
BRAM[1094]<= 32'h20A3FD09;
BRAM[1095]<= 32'hFD06F7FF;
BRAM[1096]<= 32'hF7FF2012;
BRAM[1097]<= 32'h2002FD03;
BRAM[1098]<= 32'hFD00F7FF;
BRAM[1099]<= 32'hF7FF20B2;
BRAM[1100]<= 32'h2012FCFD;
BRAM[1101]<= 32'hFCFAF7FF;
BRAM[1102]<= 32'hF7FF20FF;
BRAM[1103]<= 32'h2010FCF7;
BRAM[1104]<= 32'hFCF4F7FF;
BRAM[1105]<= 32'hF7FF2000;
BRAM[1106]<= 32'h20F8FCF1;
BRAM[1107]<= 32'hFCF8F7FF;
BRAM[1108]<= 32'hF7FF2021;
BRAM[1109]<= 32'h2004FCEB;
BRAM[1110]<= 32'hFCE8F7FF;
BRAM[1111]<= 32'hF7FF2013;
BRAM[1112]<= 32'h2036FCEF;
BRAM[1113]<= 32'hFCECF7FF;
BRAM[1114]<= 32'hF7FF2078;
BRAM[1115]<= 32'h20B4FCDF;
BRAM[1116]<= 32'hFCE6F7FF;
BRAM[1117]<= 32'hF7FF2002;
BRAM[1118]<= 32'h20B6FCD9;
BRAM[1119]<= 32'hFCE0F7FF;
BRAM[1120]<= 32'hF7FF2002;
BRAM[1121]<= 32'h2022FCD3;
BRAM[1122]<= 32'hFCD0F7FF;
BRAM[1123]<= 32'hF7FF20C1;
BRAM[1124]<= 32'h2041FCD7;
BRAM[1125]<= 32'hFCCAF7FF;
BRAM[1126]<= 32'hF7FF20C5;
BRAM[1127]<= 32'h2000FCD1;
BRAM[1128]<= 32'hFCC4F7FF;
BRAM[1129]<= 32'hF7FF2018;
BRAM[1130]<= 32'h203AFCC1;
BRAM[1131]<= 32'hFCC8F7FF;
BRAM[1132]<= 32'hF7FF2066;
BRAM[1133]<= 32'h2032FCBB;
BRAM[1134]<= 32'hF93AF000;
BRAM[1135]<= 32'hF7FF20E0;
BRAM[1136]<= 32'h200FFCBF;
BRAM[1137]<= 32'hFCB2F7FF;
BRAM[1138]<= 32'hF7FF201F;
BRAM[1139]<= 32'h201CFCAF;
BRAM[1140]<= 32'hFCACF7FF;
BRAM[1141]<= 32'hF7FF200C;
BRAM[1142]<= 32'h200FFCA9;
BRAM[1143]<= 32'hFCA6F7FF;
BRAM[1144]<= 32'hF7FF2008;
BRAM[1145]<= 32'h2048FCA3;
BRAM[1146]<= 32'hFCA0F7FF;
BRAM[1147]<= 32'hF7FF2098;
BRAM[1148]<= 32'h2037FC9D;
BRAM[1149]<= 32'hFC9AF7FF;
BRAM[1150]<= 32'hF7FF200A;
BRAM[1151]<= 32'h2013FC97;
BRAM[1152]<= 32'hFC94F7FF;
BRAM[1153]<= 32'hF7FF2004;
BRAM[1154]<= 32'h2011FC91;
BRAM[1155]<= 32'hFC8EF7FF;
BRAM[1156]<= 32'hF7FF200D;
BRAM[1157]<= 32'h2000FC8B;
BRAM[1158]<= 32'hFC88F7FF;
BRAM[1159]<= 32'hF7FF20E1;
BRAM[1160]<= 32'h200FFC8F;
BRAM[1161]<= 32'hFC82F7FF;
BRAM[1162]<= 32'hF7FF2032;
BRAM[1163]<= 32'h202EFC7F;
BRAM[1164]<= 32'hFC7CF7FF;
BRAM[1165]<= 32'hF7FF200B;
BRAM[1166]<= 32'h200DFC79;
BRAM[1167]<= 32'hFC76F7FF;
BRAM[1168]<= 32'hF7FF2005;
BRAM[1169]<= 32'h2047FC73;
BRAM[1170]<= 32'hFC70F7FF;
BRAM[1171]<= 32'hF7FF2075;
BRAM[1172]<= 32'h2037FC6D;
BRAM[1173]<= 32'hFC6AF7FF;
BRAM[1174]<= 32'hF7FF2006;
BRAM[1175]<= 32'h2010FC67;
BRAM[1176]<= 32'hFC64F7FF;
BRAM[1177]<= 32'hF7FF2003;
BRAM[1178]<= 32'h2024FC61;
BRAM[1179]<= 32'hFC5EF7FF;
BRAM[1180]<= 32'hF7FF2020;
BRAM[1181]<= 32'h2000FC5B;
BRAM[1182]<= 32'hFC58F7FF;
BRAM[1183]<= 32'hF7FF2011;
BRAM[1184]<= 32'h2078FC5F;
BRAM[1185]<= 32'hF8D4F000;
BRAM[1186]<= 32'hF7FF2029;
BRAM[1187]<= 32'h202CFC59;
BRAM[1188]<= 32'hFC56F7FF;
BRAM[1189]<= 32'h461A2300;
BRAM[1190]<= 32'h46184619;
BRAM[1191]<= 32'hF9D8F7FF;
BRAM[1192]<= 32'h4770BD10;
BRAM[1193]<= 32'h00004770;
BRAM[1194]<= 32'h2100B570;
BRAM[1195]<= 32'h220F2300;
BRAM[1196]<= 32'hB30478C4;
BRAM[1197]<= 32'h68244C15;
BRAM[1198]<= 32'h64E0F404;
BRAM[1199]<= 32'h64E0F5C4;
BRAM[1200]<= 32'hF1C10A21;
BRAM[1201]<= 32'h40CA0304;
BRAM[1202]<= 32'hFA047844;
BRAM[1203]<= 32'h7884F103;
BRAM[1204]<= 32'h43214014;
BRAM[1205]<= 32'h4C0E0109;
BRAM[1206]<= 32'h55A17806;
BRAM[1207]<= 32'hF0047804;
BRAM[1208]<= 32'h2401051F;
BRAM[1209]<= 32'h780540AC;
BRAM[1210]<= 32'h00AD116D;
BRAM[1211]<= 32'h25E0F105;
BRAM[1212]<= 32'h4100F8C5;
BRAM[1213]<= 32'h7804E009;
BRAM[1214]<= 32'h051FF004;
BRAM[1215]<= 32'h40AC2401;
BRAM[1216]<= 32'h78064D04;
BRAM[1217]<= 32'hF8451176;
BRAM[1218]<= 32'hBD704026;
BRAM[1219]<= 32'hE000ED0C;
BRAM[1220]<= 32'hE000E400;
BRAM[1221]<= 32'hE000E180;
BRAM[1222]<= 32'h43014902;
BRAM[1223]<= 32'h60114A02;
BRAM[1224]<= 32'h00004770;
BRAM[1225]<= 32'h05FA0000;
BRAM[1226]<= 32'hE000ED0C;
BRAM[1227]<= 32'h47704770;
BRAM[1228]<= 32'hB9214601;
BRAM[1229]<= 32'h69004810;
BRAM[1230]<= 32'h000FF000;
BRAM[1231]<= 32'h29014770;
BRAM[1232]<= 32'h480DD104;
BRAM[1233]<= 32'hF3C06900;
BRAM[1234]<= 32'hE7F72007;
BRAM[1235]<= 32'hD1042902;
BRAM[1236]<= 32'h69004809;
BRAM[1237]<= 32'h4007F3C0;
BRAM[1238]<= 32'h2903E7F0;
BRAM[1239]<= 32'h4806D103;
BRAM[1240]<= 32'h0E006900;
BRAM[1241]<= 32'h2904E7EA;
BRAM[1242]<= 32'h4803D103;
BRAM[1243]<= 32'hB2C06940;
BRAM[1244]<= 32'hBF00E7E4;
BRAM[1245]<= 32'h0000E7E2;
BRAM[1246]<= 32'h40001000;
BRAM[1247]<= 32'h49064805;
BRAM[1248]<= 32'h1D006048;
BRAM[1249]<= 32'h48056088;
BRAM[1250]<= 32'h01C060C8;
BRAM[1251]<= 32'h20026108;
BRAM[1252]<= 32'h47706148;
BRAM[1253]<= 32'hC0A80202;
BRAM[1254]<= 32'h40001000;
BRAM[1255]<= 32'h1F900000;
BRAM[1256]<= 32'h68004803;
BRAM[1257]<= 32'h0001F040;
BRAM[1258]<= 32'h60084901;
BRAM[1259]<= 32'h00004770;
BRAM[1260]<= 32'h40001000;
BRAM[1261]<= 32'h68004803;
BRAM[1262]<= 32'h0002F040;
BRAM[1263]<= 32'h60084901;
BRAM[1264]<= 32'h00004770;
BRAM[1265]<= 32'h40001000;
BRAM[1266]<= 32'h00004770;
BRAM[1267]<= 32'h480AB51F;
BRAM[1268]<= 32'h6008490A;
BRAM[1269]<= 32'h68004608;
BRAM[1270]<= 32'h31E1F44F;
BRAM[1271]<= 32'hF4F1FBB0;
BRAM[1272]<= 32'h90002001;
BRAM[1273]<= 32'h90029001;
BRAM[1274]<= 32'h46024603;
BRAM[1275]<= 32'h90034621;
BRAM[1276]<= 32'hF0000780;
BRAM[1277]<= 32'hBD1FFBDB;
BRAM[1278]<= 32'h02FAF080;
BRAM[1279]<= 32'h20000018;
BRAM[1280]<= 32'h47704770;
BRAM[1281]<= 32'h47704770;
BRAM[1282]<= 32'hE7FEBF00;
BRAM[1283]<= 32'h22FF21FF;
BRAM[1284]<= 32'hE006E00B;
BRAM[1285]<= 32'h1E53E001;
BRAM[1286]<= 32'h2A00B2DA;
BRAM[1287]<= 32'h1E4BDCFB;
BRAM[1288]<= 32'h2900B2D9;
BRAM[1289]<= 32'h1E43DCF6;
BRAM[1290]<= 32'h2800B2D8;
BRAM[1291]<= 32'h4770DCF1;
BRAM[1292]<= 32'h4604B510;
BRAM[1293]<= 32'h20FFE003;
BRAM[1294]<= 32'hFFE8F7FF;
BRAM[1295]<= 32'h2C001E64;
BRAM[1296]<= 32'hBD10D1F9;
BRAM[1297]<= 32'hF04F4601;
BRAM[1298]<= 32'h477030FF;
BRAM[1299]<= 32'h4604B570;
BRAM[1300]<= 32'h2C0A460D;
BRAM[1301]<= 32'h210DD103;
BRAM[1302]<= 32'hF0000740;
BRAM[1303]<= 32'h4621FB9D;
BRAM[1304]<= 32'h4080F04F;
BRAM[1305]<= 32'hFB98F000;
BRAM[1306]<= 32'hBD704620;
BRAM[1307]<= 32'h20FFB508;
BRAM[1308]<= 32'h700849FE;
BRAM[1309]<= 32'h49FE2001;
BRAM[1310]<= 32'h20007008;
BRAM[1311]<= 32'h700849FD;
BRAM[1312]<= 32'h714849FD;
BRAM[1313]<= 32'h60A0F44F;
BRAM[1314]<= 32'hFF46F7FF;
BRAM[1315]<= 32'hFEFAF7FE;
BRAM[1316]<= 32'hF8A0F7FF;
BRAM[1317]<= 32'hFE22F7FF;
BRAM[1318]<= 32'hF7FF48F8;
BRAM[1319]<= 32'h2300F906;
BRAM[1320]<= 32'h213C461A;
BRAM[1321]<= 32'hF7FF2032;
BRAM[1322]<= 32'hF44FF9E7;
BRAM[1323]<= 32'hF44F007C;
BRAM[1324]<= 32'hF44F739B;
BRAM[1325]<= 32'h213C72EB;
BRAM[1326]<= 32'hF44F9000;
BRAM[1327]<= 32'hF7FF708C;
BRAM[1328]<= 32'h2000F96F;
BRAM[1329]<= 32'h46022318;
BRAM[1330]<= 32'h90002146;
BRAM[1331]<= 32'h1023F240;
BRAM[1332]<= 32'hF98CF7FF;
BRAM[1333]<= 32'hFBCAF7FF;
BRAM[1334]<= 32'hFF50F7FF;
BRAM[1335]<= 32'hFF60F7FF;
BRAM[1336]<= 32'hF7FF200A;
BRAM[1337]<= 32'hE34DFFA5;
BRAM[1338]<= 32'h780048E2;
BRAM[1339]<= 32'h1DA1B9A8;
BRAM[1340]<= 32'h2100B2C8;
BRAM[1341]<= 32'hF889F7FF;
BRAM[1342]<= 32'hF7FF20C8;
BRAM[1343]<= 32'h1DA1FF99;
BRAM[1344]<= 32'h2101B2C8;
BRAM[1345]<= 32'hF881F7FF;
BRAM[1346]<= 32'hF7FF20C8;
BRAM[1347]<= 32'h1C60FF91;
BRAM[1348]<= 32'h2C06B2C4;
BRAM[1349]<= 32'h2400DB37;
BRAM[1350]<= 32'h48D6E035;
BRAM[1351]<= 32'h28017800;
BRAM[1352]<= 32'h1DA1D115;
BRAM[1353]<= 32'h2100B2C8;
BRAM[1354]<= 32'hF86FF7FF;
BRAM[1355]<= 32'hF7FF20C8;
BRAM[1356]<= 32'h1DA1FF7F;
BRAM[1357]<= 32'h2101B2C8;
BRAM[1358]<= 32'hF867F7FF;
BRAM[1359]<= 32'hF7FF20C8;
BRAM[1360]<= 32'h1E60FF77;
BRAM[1361]<= 32'h2C00B2C4;
BRAM[1362]<= 32'h2405DC1D;
BRAM[1363]<= 32'h48C9E01B;
BRAM[1364]<= 32'h28027800;
BRAM[1365]<= 32'hF04FD117;
BRAM[1366]<= 32'h684040A0;
BRAM[1367]<= 32'h6078F420;
BRAM[1368]<= 32'h41A0F04F;
BRAM[1369]<= 32'hF44F6048;
BRAM[1370]<= 32'hF7FF70C8;
BRAM[1371]<= 32'hF04FFF61;
BRAM[1372]<= 32'h684040A0;
BRAM[1373]<= 32'h6078F440;
BRAM[1374]<= 32'h41A0F04F;
BRAM[1375]<= 32'hF44F6048;
BRAM[1376]<= 32'hF7FF70C8;
BRAM[1377]<= 32'h48B9FF55;
BRAM[1378]<= 32'h28037800;
BRAM[1379]<= 32'h48BCD17E;
BRAM[1380]<= 32'hB2C56900;
BRAM[1381]<= 32'h23FCB93D;
BRAM[1382]<= 32'h2178A2BA;
BRAM[1383]<= 32'h70C1F44F;
BRAM[1384]<= 32'hFA2EF7FF;
BRAM[1385]<= 32'h2D02E026;
BRAM[1386]<= 32'h23FCD107;
BRAM[1387]<= 32'h2178A2B8;
BRAM[1388]<= 32'h70C1F44F;
BRAM[1389]<= 32'hFA24F7FF;
BRAM[1390]<= 32'h2D04E01C;
BRAM[1391]<= 32'h23FCD107;
BRAM[1392]<= 32'h2178A2B6;
BRAM[1393]<= 32'h70C1F44F;
BRAM[1394]<= 32'hFA1AF7FF;
BRAM[1395]<= 32'h2D05E012;
BRAM[1396]<= 32'h23FCD107;
BRAM[1397]<= 32'h2178A2B4;
BRAM[1398]<= 32'h70C1F44F;
BRAM[1399]<= 32'hFA10F7FF;
BRAM[1400]<= 32'h2D03E008;
BRAM[1401]<= 32'h23FCD106;
BRAM[1402]<= 32'h2178A2AF;
BRAM[1403]<= 32'h70C1F44F;
BRAM[1404]<= 32'hFA06F7FF;
BRAM[1405]<= 32'h698048A2;
BRAM[1406]<= 32'h2015F3C0;
BRAM[1407]<= 32'h600849AD;
BRAM[1408]<= 32'h68004608;
BRAM[1409]<= 32'h7110F242;
BRAM[1410]<= 32'hF0F1FBB0;
BRAM[1411]<= 32'h499A3030;
BRAM[1412]<= 32'h48A87008;
BRAM[1413]<= 32'hF2426800;
BRAM[1414]<= 32'hFBB07110;
BRAM[1415]<= 32'hFB01F2F1;
BRAM[1416]<= 32'hF44F0012;
BRAM[1417]<= 32'hFBB0717A;
BRAM[1418]<= 32'h3030F0F1;
BRAM[1419]<= 32'h70484992;
BRAM[1420]<= 32'h680048A0;
BRAM[1421]<= 32'h7110F242;
BRAM[1422]<= 32'hF2F1FBB0;
BRAM[1423]<= 32'h0012FB01;
BRAM[1424]<= 32'h717AF44F;
BRAM[1425]<= 32'hF2F1FBB0;
BRAM[1426]<= 32'h0012FB01;
BRAM[1427]<= 32'hFBB02164;
BRAM[1428]<= 32'h3030F0F1;
BRAM[1429]<= 32'h70884988;
BRAM[1430]<= 32'h68004896;
BRAM[1431]<= 32'h7110F242;
BRAM[1432]<= 32'hF2F1FBB0;
BRAM[1433]<= 32'h0012FB01;
BRAM[1434]<= 32'h717AF44F;
BRAM[1435]<= 32'hF2F1FBB0;
BRAM[1436]<= 32'h0012FB01;
BRAM[1437]<= 32'hFBB02164;
BRAM[1438]<= 32'hFB01F2F1;
BRAM[1439]<= 32'h210A0012;
BRAM[1440]<= 32'hF0F1FBB0;
BRAM[1441]<= 32'h497C3030;
BRAM[1442]<= 32'hE00070C8;
BRAM[1443]<= 32'h4889E271;
BRAM[1444]<= 32'hF2426800;
BRAM[1445]<= 32'hFBB07110;
BRAM[1446]<= 32'hFB01F2F1;
BRAM[1447]<= 32'hF44F0012;
BRAM[1448]<= 32'hFBB0717A;
BRAM[1449]<= 32'hFB01F2F1;
BRAM[1450]<= 32'h21640012;
BRAM[1451]<= 32'hF2F1FBB0;
BRAM[1452]<= 32'h0012FB01;
BRAM[1453]<= 32'hFBB0210A;
BRAM[1454]<= 32'hFB01F2F1;
BRAM[1455]<= 32'h30300012;
BRAM[1456]<= 32'h7108496D;
BRAM[1457]<= 32'h71482000;
BRAM[1458]<= 32'h460A23FC;
BRAM[1459]<= 32'hF44F2190;
BRAM[1460]<= 32'hF7FF70C1;
BRAM[1461]<= 32'h486AF995;
BRAM[1462]<= 32'hF3C069C0;
BRAM[1463]<= 32'h497510D5;
BRAM[1464]<= 32'h46086008;
BRAM[1465]<= 32'hF2426800;
BRAM[1466]<= 32'hFBB07110;
BRAM[1467]<= 32'h3030F0F1;
BRAM[1468]<= 32'h70084961;
BRAM[1469]<= 32'h6800486F;
BRAM[1470]<= 32'h7110F242;
BRAM[1471]<= 32'hF2F1FBB0;
BRAM[1472]<= 32'h0012FB01;
BRAM[1473]<= 32'h717AF44F;
BRAM[1474]<= 32'hF0F1FBB0;
BRAM[1475]<= 32'h495A3030;
BRAM[1476]<= 32'h48687048;
BRAM[1477]<= 32'hF2426800;
BRAM[1478]<= 32'hFBB07110;
BRAM[1479]<= 32'hFB01F2F1;
BRAM[1480]<= 32'hF44F0012;
BRAM[1481]<= 32'hFBB0717A;
BRAM[1482]<= 32'hFB01F2F1;
BRAM[1483]<= 32'h21640012;
BRAM[1484]<= 32'hF0F1FBB0;
BRAM[1485]<= 32'h49503030;
BRAM[1486]<= 32'h485E7088;
BRAM[1487]<= 32'hF2426800;
BRAM[1488]<= 32'hFBB07110;
BRAM[1489]<= 32'hFB01F2F1;
BRAM[1490]<= 32'hF44F0012;
BRAM[1491]<= 32'hFBB0717A;
BRAM[1492]<= 32'hFB01F2F1;
BRAM[1493]<= 32'h21640012;
BRAM[1494]<= 32'hF2F1FBB0;
BRAM[1495]<= 32'h0012FB01;
BRAM[1496]<= 32'hFBB0210A;
BRAM[1497]<= 32'h3030F0F1;
BRAM[1498]<= 32'h70C84943;
BRAM[1499]<= 32'h68004851;
BRAM[1500]<= 32'h7110F242;
BRAM[1501]<= 32'hF2F1FBB0;
BRAM[1502]<= 32'h0012FB01;
BRAM[1503]<= 32'h717AF44F;
BRAM[1504]<= 32'hF2F1FBB0;
BRAM[1505]<= 32'h0012FB01;
BRAM[1506]<= 32'hFBB02164;
BRAM[1507]<= 32'hFB01F2F1;
BRAM[1508]<= 32'h210A0012;
BRAM[1509]<= 32'hF2F1FBB0;
BRAM[1510]<= 32'h0012FB01;
BRAM[1511]<= 32'h49363030;
BRAM[1512]<= 32'h20007108;
BRAM[1513]<= 32'h23FC7148;
BRAM[1514]<= 32'h21A8460A;
BRAM[1515]<= 32'h70C1F44F;
BRAM[1516]<= 32'hF926F7FF;
BRAM[1517]<= 32'h6A004832;
BRAM[1518]<= 32'h493EB2C0;
BRAM[1519]<= 32'h46086008;
BRAM[1520]<= 32'h21646800;
BRAM[1521]<= 32'hF0F1FBB0;
BRAM[1522]<= 32'h492B3030;
BRAM[1523]<= 32'h48397008;
BRAM[1524]<= 32'h21646800;
BRAM[1525]<= 32'hF2F1FBB0;
BRAM[1526]<= 32'h0012FB01;
BRAM[1527]<= 32'hFBB0210A;
BRAM[1528]<= 32'h3030F0F1;
BRAM[1529]<= 32'h70484924;
BRAM[1530]<= 32'h68004832;
BRAM[1531]<= 32'hFBB02164;
BRAM[1532]<= 32'hFB01F2F1;
BRAM[1533]<= 32'h210A0012;
BRAM[1534]<= 32'hF2F1FBB0;
BRAM[1535]<= 32'h0012FB01;
BRAM[1536]<= 32'h491D3030;
BRAM[1537]<= 32'h20007088;
BRAM[1538]<= 32'h23FC70C8;
BRAM[1539]<= 32'h21C0460A;
BRAM[1540]<= 32'h70C1F44F;
BRAM[1541]<= 32'hF8F4F7FF;
BRAM[1542]<= 32'h6A004819;
BRAM[1543]<= 32'h2007F3C0;
BRAM[1544]<= 32'h49240040;
BRAM[1545]<= 32'h46086008;
BRAM[1546]<= 32'h21646800;
BRAM[1547]<= 32'hF0F1FBB0;
BRAM[1548]<= 32'h49113030;
BRAM[1549]<= 32'h481F7008;
BRAM[1550]<= 32'h21646800;
BRAM[1551]<= 32'hF2F1FBB0;
BRAM[1552]<= 32'h0012FB01;
BRAM[1553]<= 32'hFBB0210A;
BRAM[1554]<= 32'h3030F0F1;
BRAM[1555]<= 32'h7048490A;
BRAM[1556]<= 32'h68004818;
BRAM[1557]<= 32'hFBB02164;
BRAM[1558]<= 32'hFB01F2F1;
BRAM[1559]<= 32'h210A0012;
BRAM[1560]<= 32'hF2F1FBB0;
BRAM[1561]<= 32'h0012FB01;
BRAM[1562]<= 32'hE0253030;
BRAM[1563]<= 32'h2000000D;
BRAM[1564]<= 32'h2000000E;
BRAM[1565]<= 32'h2000000C;
BRAM[1566]<= 32'h20000000;
BRAM[1567]<= 32'h00FCFCFC;
BRAM[1568]<= 32'h40001000;
BRAM[1569]<= 32'h454C4449;
BRAM[1570]<= 32'h20202020;
BRAM[1571]<= 32'h00000000;
BRAM[1572]<= 32'h646E6553;
BRAM[1573]<= 32'h4E595320;
BRAM[1574]<= 32'h00000000;
BRAM[1575]<= 32'h646E6553;
BRAM[1576]<= 32'h4B434120;
BRAM[1577]<= 32'h00000000;
BRAM[1578]<= 32'h65636552;
BRAM[1579]<= 32'h20657669;
BRAM[1580]<= 32'h00000000;
BRAM[1581]<= 32'h20000008;
BRAM[1582]<= 32'h708849B3;
BRAM[1583]<= 32'h70C82000;
BRAM[1584]<= 32'h460A23FC;
BRAM[1585]<= 32'hF44F21D8;
BRAM[1586]<= 32'hF7FF70C1;
BRAM[1587]<= 32'h48AFF899;
BRAM[1588]<= 32'hB2806A40;
BRAM[1589]<= 32'h600849AE;
BRAM[1590]<= 32'h68004608;
BRAM[1591]<= 32'h7110F242;
BRAM[1592]<= 32'hF0F1FBB0;
BRAM[1593]<= 32'h49A83030;
BRAM[1594]<= 32'h48A97008;
BRAM[1595]<= 32'hF2426800;
BRAM[1596]<= 32'hFBB07110;
BRAM[1597]<= 32'hFB01F2F1;
BRAM[1598]<= 32'hF44F0012;
BRAM[1599]<= 32'hFBB0717A;
BRAM[1600]<= 32'h3030F0F1;
BRAM[1601]<= 32'h704849A0;
BRAM[1602]<= 32'h680048A1;
BRAM[1603]<= 32'h7110F242;
BRAM[1604]<= 32'hF2F1FBB0;
BRAM[1605]<= 32'h0012FB01;
BRAM[1606]<= 32'h717AF44F;
BRAM[1607]<= 32'hF2F1FBB0;
BRAM[1608]<= 32'h0012FB01;
BRAM[1609]<= 32'hFBB02164;
BRAM[1610]<= 32'h3030F0F1;
BRAM[1611]<= 32'h70884996;
BRAM[1612]<= 32'h68004897;
BRAM[1613]<= 32'h7110F242;
BRAM[1614]<= 32'hF2F1FBB0;
BRAM[1615]<= 32'h0012FB01;
BRAM[1616]<= 32'h717AF44F;
BRAM[1617]<= 32'hF2F1FBB0;
BRAM[1618]<= 32'h0012FB01;
BRAM[1619]<= 32'hFBB02164;
BRAM[1620]<= 32'hFB01F2F1;
BRAM[1621]<= 32'h210A0012;
BRAM[1622]<= 32'hF0F1FBB0;
BRAM[1623]<= 32'h498A3030;
BRAM[1624]<= 32'h488B70C8;
BRAM[1625]<= 32'hF2426800;
BRAM[1626]<= 32'hFBB07110;
BRAM[1627]<= 32'hFB01F2F1;
BRAM[1628]<= 32'hF44F0012;
BRAM[1629]<= 32'hFBB0717A;
BRAM[1630]<= 32'hFB01F2F1;
BRAM[1631]<= 32'h21640012;
BRAM[1632]<= 32'hF2F1FBB0;
BRAM[1633]<= 32'h0012FB01;
BRAM[1634]<= 32'hFBB0210A;
BRAM[1635]<= 32'hFB01F2F1;
BRAM[1636]<= 32'h30300012;
BRAM[1637]<= 32'h7108497C;
BRAM[1638]<= 32'h71482000;
BRAM[1639]<= 32'h460A23FC;
BRAM[1640]<= 32'hF44F21F0;
BRAM[1641]<= 32'hF7FF70C1;
BRAM[1642]<= 32'h4878F82B;
BRAM[1643]<= 32'hF64F6A40;
BRAM[1644]<= 32'hEA0171FF;
BRAM[1645]<= 32'h49764010;
BRAM[1646]<= 32'h46086008;
BRAM[1647]<= 32'hF2426800;
BRAM[1648]<= 32'hFBB07110;
BRAM[1649]<= 32'h3030F0F1;
BRAM[1650]<= 32'h7008496F;
BRAM[1651]<= 32'h68004870;
BRAM[1652]<= 32'h7110F242;
BRAM[1653]<= 32'hF2F1FBB0;
BRAM[1654]<= 32'h0012FB01;
BRAM[1655]<= 32'h717AF44F;
BRAM[1656]<= 32'hF0F1FBB0;
BRAM[1657]<= 32'h49683030;
BRAM[1658]<= 32'h48697048;
BRAM[1659]<= 32'hF2426800;
BRAM[1660]<= 32'hFBB07110;
BRAM[1661]<= 32'hFB01F2F1;
BRAM[1662]<= 32'hF44F0012;
BRAM[1663]<= 32'hFBB0717A;
BRAM[1664]<= 32'hFB01F2F1;
BRAM[1665]<= 32'h21640012;
BRAM[1666]<= 32'hF0F1FBB0;
BRAM[1667]<= 32'h495E3030;
BRAM[1668]<= 32'h485F7088;
BRAM[1669]<= 32'hF2426800;
BRAM[1670]<= 32'hFBB07110;
BRAM[1671]<= 32'hFB01F2F1;
BRAM[1672]<= 32'hF44F0012;
BRAM[1673]<= 32'hFBB0717A;
BRAM[1674]<= 32'hFB01F2F1;
BRAM[1675]<= 32'h21640012;
BRAM[1676]<= 32'hF2F1FBB0;
BRAM[1677]<= 32'h0012FB01;
BRAM[1678]<= 32'hFBB0210A;
BRAM[1679]<= 32'h3030F0F1;
BRAM[1680]<= 32'h70C84951;
BRAM[1681]<= 32'h68004852;
BRAM[1682]<= 32'h7110F242;
BRAM[1683]<= 32'hF2F1FBB0;
BRAM[1684]<= 32'h0012FB01;
BRAM[1685]<= 32'h717AF44F;
BRAM[1686]<= 32'hF2F1FBB0;
BRAM[1687]<= 32'h0012FB01;
BRAM[1688]<= 32'hFBB02164;
BRAM[1689]<= 32'hFB01F2F1;
BRAM[1690]<= 32'h210A0012;
BRAM[1691]<= 32'hF2F1FBB0;
BRAM[1692]<= 32'h0012FB01;
BRAM[1693]<= 32'h49443030;
BRAM[1694]<= 32'h20007108;
BRAM[1695]<= 32'h23FC7148;
BRAM[1696]<= 32'hF44F460A;
BRAM[1697]<= 32'hF44F7184;
BRAM[1698]<= 32'hF7FE70C1;
BRAM[1699]<= 32'h483FFFB9;
BRAM[1700]<= 32'hF64F6A00;
BRAM[1701]<= 32'hEA0171FF;
BRAM[1702]<= 32'h493D4010;
BRAM[1703]<= 32'h46086008;
BRAM[1704]<= 32'hF2426800;
BRAM[1705]<= 32'hFBB07110;
BRAM[1706]<= 32'h3030F0F1;
BRAM[1707]<= 32'h70084936;
BRAM[1708]<= 32'h68004837;
BRAM[1709]<= 32'h7110F242;
BRAM[1710]<= 32'hF2F1FBB0;
BRAM[1711]<= 32'h0012FB01;
BRAM[1712]<= 32'h717AF44F;
BRAM[1713]<= 32'hF0F1FBB0;
BRAM[1714]<= 32'h492F3030;
BRAM[1715]<= 32'h48307048;
BRAM[1716]<= 32'hF2426800;
BRAM[1717]<= 32'hFBB07110;
BRAM[1718]<= 32'hFB01F2F1;
BRAM[1719]<= 32'hF44F0012;
BRAM[1720]<= 32'hFBB0717A;
BRAM[1721]<= 32'hFB01F2F1;
BRAM[1722]<= 32'h21640012;
BRAM[1723]<= 32'hF0F1FBB0;
BRAM[1724]<= 32'h49253030;
BRAM[1725]<= 32'h48267088;
BRAM[1726]<= 32'hF2426800;
BRAM[1727]<= 32'hFBB07110;
BRAM[1728]<= 32'hFB01F2F1;
BRAM[1729]<= 32'hF44F0012;
BRAM[1730]<= 32'hFBB0717A;
BRAM[1731]<= 32'hFB01F2F1;
BRAM[1732]<= 32'h21640012;
BRAM[1733]<= 32'hF2F1FBB0;
BRAM[1734]<= 32'h0012FB01;
BRAM[1735]<= 32'hFBB0210A;
BRAM[1736]<= 32'h3030F0F1;
BRAM[1737]<= 32'h70C84918;
BRAM[1738]<= 32'h68004819;
BRAM[1739]<= 32'h7110F242;
BRAM[1740]<= 32'hF2F1FBB0;
BRAM[1741]<= 32'h0012FB01;
BRAM[1742]<= 32'h717AF44F;
BRAM[1743]<= 32'hF2F1FBB0;
BRAM[1744]<= 32'h0012FB01;
BRAM[1745]<= 32'hFBB02164;
BRAM[1746]<= 32'hFB01F2F1;
BRAM[1747]<= 32'h210A0012;
BRAM[1748]<= 32'hF2F1FBB0;
BRAM[1749]<= 32'h0012FB01;
BRAM[1750]<= 32'h490B3030;
BRAM[1751]<= 32'h20007108;
BRAM[1752]<= 32'h23FC7148;
BRAM[1753]<= 32'hF44F460A;
BRAM[1754]<= 32'hF44F7190;
BRAM[1755]<= 32'hF7FE70C1;
BRAM[1756]<= 32'h4808FF47;
BRAM[1757]<= 32'h28017800;
BRAM[1758]<= 32'h2000D104;
BRAM[1759]<= 32'h70084905;
BRAM[1760]<= 32'hF874F7FF;
BRAM[1761]<= 32'h0000E4B0;
BRAM[1762]<= 32'h20000000;
BRAM[1763]<= 32'h40001000;
BRAM[1764]<= 32'h20000008;
BRAM[1765]<= 32'h2000000F;
BRAM[1766]<= 32'h6842E004;
BRAM[1767]<= 32'h0201F002;
BRAM[1768]<= 32'hE000B902;
BRAM[1769]<= 32'hBF00E7F9;
BRAM[1770]<= 32'h47706001;
BRAM[1771]<= 32'h41F0E92D;
BRAM[1772]<= 32'h460D4604;
BRAM[1773]<= 32'hC808E9DD;
BRAM[1774]<= 32'h6706E9DD;
BRAM[1775]<= 32'hB10A2100;
BRAM[1776]<= 32'h0101F041;
BRAM[1777]<= 32'hF041B10B;
BRAM[1778]<= 32'hB10E0102;
BRAM[1779]<= 32'h0104F041;
BRAM[1780]<= 32'hF041B10F;
BRAM[1781]<= 32'hF1BC0108;
BRAM[1782]<= 32'hD0010F00;
BRAM[1783]<= 32'h0110F041;
BRAM[1784]<= 32'h0F00F1B8;
BRAM[1785]<= 32'hF041D001;
BRAM[1786]<= 32'h20000120;
BRAM[1787]<= 32'h612560A0;
BRAM[1788]<= 32'h686060A1;
BRAM[1789]<= 32'h000CF000;
BRAM[1790]<= 32'h2001B110;
BRAM[1791]<= 32'h81F0E8BD;
BRAM[1792]<= 32'hE7FB2000;
BRAM[1793]<= 32'h00000000;
BRAM[1794]<= 32'h00000000;
BRAM[1795]<= 32'h00000000;
BRAM[1796]<= 32'h80000180;
BRAM[1797]<= 32'hD9800001;
BRAM[1798]<= 32'h0FDFE00C;
BRAM[1799]<= 32'h800CD980;
BRAM[1800]<= 32'hD9800CD9;
BRAM[1801]<= 32'h0CD9800C;
BRAM[1802]<= 32'h800CD980;
BRAM[1803]<= 32'hD9800CD9;
BRAM[1804]<= 32'h0CD9800C;
BRAM[1805]<= 32'h800CD980;
BRAM[1806]<= 32'hD9800CD9;
BRAM[1807]<= 32'h0CD9800C;
BRAM[1808]<= 32'h400CD880;
BRAM[1809]<= 32'hCE200FD8;
BRAM[1810]<= 32'h0001100C;
BRAM[1811]<= 32'h00000000;
BRAM[1812]<= 32'h00000000;
BRAM[1813]<= 32'h00000000;
BRAM[1814]<= 32'h40006000;
BRAM[1815]<= 32'hFCC00060;
BRAM[1816]<= 32'h00608007;
BRAM[1817]<= 32'h00066480;
BRAM[1818]<= 32'h64F007FC;
BRAM[1819]<= 32'h0664C006;
BRAM[1820]<= 32'hC007FCC0;
BRAM[1821]<= 32'hF0C006E4;
BRAM[1822]<= 32'h0170C000;
BRAM[1823]<= 32'hC00378C0;
BRAM[1824]<= 32'h64C00668;
BRAM[1825]<= 32'h0462C006;
BRAM[1826]<= 32'h700060C0;
BRAM[1827]<= 32'hFE300001;
BRAM[1828]<= 32'h00000007;
BRAM[1829]<= 32'h00000000;
BRAM[1830]<= 32'h00000000;
BRAM[1831]<= 32'h06000000;
BRAM[1832]<= 32'hC007EFC0;
BRAM[1833]<= 32'h6CC0066C;
BRAM[1834]<= 32'h066CC006;
BRAM[1835]<= 32'hC0066CC0;
BRAM[1836]<= 32'h90C007EF;
BRAM[1837]<= 32'h01180000;
BRAM[1838]<= 32'h000FFFE0;
BRAM[1839]<= 32'h8200004C;
BRAM[1840]<= 32'h1F018001;
BRAM[1841]<= 32'hC01FEFE0;
BRAM[1842]<= 32'h6CC0066C;
BRAM[1843]<= 32'h066CC006;
BRAM[1844]<= 32'hC0066CC0;
BRAM[1845]<= 32'h6CC007EF;
BRAM[1846]<= 32'h00000006;
BRAM[1847]<= 32'h00000000;
BRAM[1848]<= 32'h00000000;
BRAM[1849]<= 32'h00C30000;
BRAM[1850]<= 32'h0000C300;
BRAM[1851]<= 32'hC30001C3;
BRAM[1852]<= 32'h06C31002;
BRAM[1853]<= 32'h2004C320;
BRAM[1854]<= 32'hFF6000C3;
BRAM[1855]<= 32'h00C3000F;
BRAM[1856]<= 32'h0000C300;
BRAM[1857]<= 32'hC38000C3;
BRAM[1858]<= 32'h00C34000;
BRAM[1859]<= 32'h3000E370;
BRAM[1860]<= 32'h23100163;
BRAM[1861]<= 32'h07330003;
BRAM[1862]<= 32'h000E1300;
BRAM[1863]<= 32'h07000C0B;
BRAM[1864]<= 32'h0004000C;
BRAM[1865]<= 32'h00000000;
BRAM[1866]<= 32'h00000000;
BRAM[1867]<= 32'h00000000;
BRAM[1868]<= 32'h00001800;
BRAM[1869]<= 32'h18000018;
BRAM[1870]<= 32'h0FFFE000;
BRAM[1871]<= 32'h00003800;
BRAM[1872]<= 32'h84000048;
BRAM[1873]<= 32'h018A0000;
BRAM[1874]<= 32'h800F3100;
BRAM[1875]<= 32'h20600C20;
BRAM[1876]<= 32'h0016C008;
BRAM[1877]<= 32'hC00226C0;
BRAM[1878]<= 32'h66C00666;
BRAM[1879]<= 32'h0D06C005;
BRAM[1880]<= 32'h400906C0;
BRAM[1881]<= 32'hFE200106;
BRAM[1882]<= 32'h00000001;
BRAM[1883]<= 32'h00000000;
BRAM[1884]<= 32'h00000000;
BRAM[1885]<= 32'h00040000;
BRAM[1886]<= 32'hC000C4C0;
BRAM[1887]<= 32'hC4C000C4;
BRAM[1888]<= 32'h0044C00F;
BRAM[1889]<= 32'hC00064C0;
BRAM[1890]<= 32'h14C000A4;
BRAM[1891]<= 32'h0304C001;
BRAM[1892]<= 32'h000204C0;
BRAM[1893]<= 32'h00000204;
BRAM[1894]<= 32'h03FFC000;
BRAM[1895]<= 32'hC00364C0;
BRAM[1896]<= 32'h64C00364;
BRAM[1897]<= 32'h0364C003;
BRAM[1898]<= 32'hC00364C0;
BRAM[1899]<= 32'hFFF00364;
BRAM[1900]<= 32'h0000000F;
BRAM[1901]<= 32'h00000000;
BRAM[1902]<= 32'h00000000;
BRAM[1903]<= 32'h00000000;
BRAM[1904]<= 32'h8000C180;
BRAM[1905]<= 32'hFD800081;
BRAM[1906]<= 32'h0C0D800F;
BRAM[1907]<= 32'h80040FF0;
BRAM[1908]<= 32'h21800361;
BRAM[1909]<= 32'h06358002;
BRAM[1910]<= 32'hC00C1380;
BRAM[1911]<= 32'h01F00C09;
BRAM[1912]<= 32'h0FF9A000;
BRAM[1913]<= 32'h8000C180;
BRAM[1914]<= 32'hC18000C1;
BRAM[1915]<= 32'h00C18000;
BRAM[1916]<= 32'h8000C180;
BRAM[1917]<= 32'hFCE000C1;
BRAM[1918]<= 32'h0000001F;
BRAM[1919]<= 32'h18000000;
BRAM[1920]<= 32'h42424224;
BRAM[1921]<= 32'h42424242;
BRAM[1922]<= 32'h00001824;
BRAM[1923]<= 32'h10000000;
BRAM[1924]<= 32'h1010101C;
BRAM[1925]<= 32'h10101010;
BRAM[1926]<= 32'h00007C10;
BRAM[1927]<= 32'h3C000000;
BRAM[1928]<= 32'h40424242;
BRAM[1929]<= 32'h04081020;
BRAM[1930]<= 32'h00007E42;
BRAM[1931]<= 32'h3C000000;
BRAM[1932]<= 32'h20404242;
BRAM[1933]<= 32'h42402018;
BRAM[1934]<= 32'h00003C42;
BRAM[1935]<= 32'h20000000;
BRAM[1936]<= 32'h24283030;
BRAM[1937]<= 32'h20FE2224;
BRAM[1938]<= 32'h0000F820;
BRAM[1939]<= 32'h7E000000;
BRAM[1940]<= 32'h1E020202;
BRAM[1941]<= 32'h42404022;
BRAM[1942]<= 32'h00001C22;
BRAM[1943]<= 32'h18000000;
BRAM[1944]<= 32'h3A020224;
BRAM[1945]<= 32'h42424246;
BRAM[1946]<= 32'h00003844;
BRAM[1947]<= 32'h7E000000;
BRAM[1948]<= 32'h10202042;
BRAM[1949]<= 32'h08080810;
BRAM[1950]<= 32'h00000808;
BRAM[1951]<= 32'h3C000000;
BRAM[1952]<= 32'h24424242;
BRAM[1953]<= 32'h42422418;
BRAM[1954]<= 32'h00003C42;
BRAM[1955]<= 32'h1C000000;
BRAM[1956]<= 32'h42424222;
BRAM[1957]<= 32'h40405C62;
BRAM[1958]<= 32'h00001824;
BRAM[1959]<= 32'h08000000;
BRAM[1960]<= 32'h14141808;
BRAM[1961]<= 32'h42223C24;
BRAM[1962]<= 32'h0000E742;
BRAM[1963]<= 32'h1F000000;
BRAM[1964]<= 32'h1E222222;
BRAM[1965]<= 32'h42424222;
BRAM[1966]<= 32'h00001F22;
BRAM[1967]<= 32'h7C000000;
BRAM[1968]<= 32'h01014242;
BRAM[1969]<= 32'h42010101;
BRAM[1970]<= 32'h00001C22;
BRAM[1971]<= 32'h1F000000;
BRAM[1972]<= 32'h42424222;
BRAM[1973]<= 32'h42424242;
BRAM[1974]<= 32'h00001F22;
BRAM[1975]<= 32'h3F000000;
BRAM[1976]<= 32'h1E121242;
BRAM[1977]<= 32'h42021212;
BRAM[1978]<= 32'h00003F42;
BRAM[1979]<= 32'h3F000000;
BRAM[1980]<= 32'h1E121242;
BRAM[1981]<= 32'h02021212;
BRAM[1982]<= 32'h00000702;
BRAM[1983]<= 32'h3C000000;
BRAM[1984]<= 32'h01012222;
BRAM[1985]<= 32'h22217101;
BRAM[1986]<= 32'h00001C22;
BRAM[1987]<= 32'hE7000000;
BRAM[1988]<= 32'h42424242;
BRAM[1989]<= 32'h4242427E;
BRAM[1990]<= 32'h0000E742;
BRAM[1991]<= 32'h3E000000;
BRAM[1992]<= 32'h08080808;
BRAM[1993]<= 32'h08080808;
BRAM[1994]<= 32'h00003E08;
BRAM[1995]<= 32'h7C000000;
BRAM[1996]<= 32'h10101010;
BRAM[1997]<= 32'h10101010;
BRAM[1998]<= 32'h0F111010;
BRAM[1999]<= 32'h77000000;
BRAM[2000]<= 32'h0E0A1222;
BRAM[2001]<= 32'h2212120A;
BRAM[2002]<= 32'h00007722;
BRAM[2003]<= 32'h07000000;
BRAM[2004]<= 32'h02020202;
BRAM[2005]<= 32'h02020202;
BRAM[2006]<= 32'h00007F42;
BRAM[2007]<= 32'h77000000;
BRAM[2008]<= 32'h36363636;
BRAM[2009]<= 32'h2A2A2A36;
BRAM[2010]<= 32'h00006B2A;
BRAM[2011]<= 32'hE3000000;
BRAM[2012]<= 32'h4A4A4646;
BRAM[2013]<= 32'h62525252;
BRAM[2014]<= 32'h00004762;
BRAM[2015]<= 32'h1C000000;
BRAM[2016]<= 32'h41414122;
BRAM[2017]<= 32'h41414141;
BRAM[2018]<= 32'h00001C22;
BRAM[2019]<= 32'h3F000000;
BRAM[2020]<= 32'h42424242;
BRAM[2021]<= 32'h0202023E;
BRAM[2022]<= 32'h00000702;
BRAM[2023]<= 32'h1C000000;
BRAM[2024]<= 32'h41414122;
BRAM[2025]<= 32'h4D414141;
BRAM[2026]<= 32'h00601C32;
BRAM[2027]<= 32'h3F000000;
BRAM[2028]<= 32'h3E424242;
BRAM[2029]<= 32'h22221212;
BRAM[2030]<= 32'h0000C742;
BRAM[2031]<= 32'h7C000000;
BRAM[2032]<= 32'h04024242;
BRAM[2033]<= 32'h42402018;
BRAM[2034]<= 32'h00003E42;
BRAM[2035]<= 32'h7F000000;
BRAM[2036]<= 32'h08080849;
BRAM[2037]<= 32'h08080808;
BRAM[2038]<= 32'h00001C08;
BRAM[2039]<= 32'hE7000000;
BRAM[2040]<= 32'h42424242;
BRAM[2041]<= 32'h42424242;
BRAM[2042]<= 32'h00003C42;
BRAM[2043]<= 32'hE7000000;
BRAM[2044]<= 32'h24224242;
BRAM[2045]<= 32'h18141424;
BRAM[2046]<= 32'h00000808;
BRAM[2047]<= 32'h6B000000;
BRAM[2048]<= 32'h2A2A2A2A;
BRAM[2049]<= 32'h1414362A;
BRAM[2050]<= 32'h00001414;
BRAM[2051]<= 32'hE7000000;
BRAM[2052]<= 32'h18242442;
BRAM[2053]<= 32'h24241818;
BRAM[2054]<= 32'h0000E742;
BRAM[2055]<= 32'h77000000;
BRAM[2056]<= 32'h14142222;
BRAM[2057]<= 32'h08080808;
BRAM[2058]<= 32'h00001C08;
BRAM[2059]<= 32'h7E000000;
BRAM[2060]<= 32'h10102021;
BRAM[2061]<= 32'h42040408;
BRAM[2062]<= 32'h00003F42;
BRAM[2063]<= 32'h00000000;
BRAM[2064]<= 32'h1C000000;
BRAM[2065]<= 32'h222C3022;
BRAM[2066]<= 32'h00006C32;
BRAM[2067]<= 32'h00000000;
BRAM[2068]<= 32'h1A020203;
BRAM[2069]<= 32'h42424226;
BRAM[2070]<= 32'h00001A26;
BRAM[2071]<= 32'h00000000;
BRAM[2072]<= 32'h38000000;
BRAM[2073]<= 32'h02020244;
BRAM[2074]<= 32'h00003844;
BRAM[2075]<= 32'h00000000;
BRAM[2076]<= 32'h7C404060;
BRAM[2077]<= 32'h42424242;
BRAM[2078]<= 32'h0000DC62;
BRAM[2079]<= 32'h00000000;
BRAM[2080]<= 32'h3C000000;
BRAM[2081]<= 32'h027E4242;
BRAM[2082]<= 32'h00003C42;
BRAM[2083]<= 32'h00000000;
BRAM[2084]<= 32'h3E084830;
BRAM[2085]<= 32'h08080808;
BRAM[2086]<= 32'h00003E08;
BRAM[2087]<= 32'h00000000;
BRAM[2088]<= 32'h7C000000;
BRAM[2089]<= 32'h021C2222;
BRAM[2090]<= 32'h3C42423C;
BRAM[2091]<= 32'h00000000;
BRAM[2092]<= 32'h3A020203;
BRAM[2093]<= 32'h42424246;
BRAM[2094]<= 32'h0000E742;
BRAM[2095]<= 32'h0C000000;
BRAM[2096]<= 32'h0E00000C;
BRAM[2097]<= 32'h08080808;
BRAM[2098]<= 32'h00003E08;
BRAM[2099]<= 32'h30000000;
BRAM[2100]<= 32'h38000030;
BRAM[2101]<= 32'h20202020;
BRAM[2102]<= 32'h1E222020;
BRAM[2103]<= 32'h00000000;
BRAM[2104]<= 32'h72020203;
BRAM[2105]<= 32'h120E0A12;
BRAM[2106]<= 32'h00007722;
BRAM[2107]<= 32'h08000000;
BRAM[2108]<= 32'h0808080E;
BRAM[2109]<= 32'h08080808;
BRAM[2110]<= 32'h00003E08;
BRAM[2111]<= 32'h00000000;
BRAM[2112]<= 32'h7F000000;
BRAM[2113]<= 32'h92929292;
BRAM[2114]<= 32'h0000B792;
BRAM[2115]<= 32'h00000000;
BRAM[2116]<= 32'h3B000000;
BRAM[2117]<= 32'h42424246;
BRAM[2118]<= 32'h0000E742;
BRAM[2119]<= 32'h00000000;
BRAM[2120]<= 32'h3C000000;
BRAM[2121]<= 32'h42424242;
BRAM[2122]<= 32'h00003C42;
BRAM[2123]<= 32'h00000000;
BRAM[2124]<= 32'h1B000000;
BRAM[2125]<= 32'h42424226;
BRAM[2126]<= 32'h07021A26;
BRAM[2127]<= 32'h00000000;
BRAM[2128]<= 32'h58000000;
BRAM[2129]<= 32'h42424264;
BRAM[2130]<= 32'hE0405864;
BRAM[2131]<= 32'h00000000;
BRAM[2132]<= 32'h77000000;
BRAM[2133]<= 32'h0404044C;
BRAM[2134]<= 32'h00001F04;
BRAM[2135]<= 32'h00000000;
BRAM[2136]<= 32'h7C000000;
BRAM[2137]<= 32'h403C0242;
BRAM[2138]<= 32'h00003E42;
BRAM[2139]<= 32'h00000000;
BRAM[2140]<= 32'h3E080800;
BRAM[2141]<= 32'h08080808;
BRAM[2142]<= 32'h00003048;
BRAM[2143]<= 32'h00000000;
BRAM[2144]<= 32'h63000000;
BRAM[2145]<= 32'h42424242;
BRAM[2146]<= 32'h0000DC62;
BRAM[2147]<= 32'h00000000;
BRAM[2148]<= 32'h77000000;
BRAM[2149]<= 32'h14142222;
BRAM[2150]<= 32'h00000808;
BRAM[2151]<= 32'h00000000;
BRAM[2152]<= 32'hDB000000;
BRAM[2153]<= 32'h2A5A5291;
BRAM[2154]<= 32'h00002424;
BRAM[2155]<= 32'h00000000;
BRAM[2156]<= 32'h6E000000;
BRAM[2157]<= 32'h18181824;
BRAM[2158]<= 32'h00007624;
BRAM[2159]<= 32'h00000000;
BRAM[2160]<= 32'hE7000000;
BRAM[2161]<= 32'h18242442;
BRAM[2162]<= 32'h06080818;
BRAM[2163]<= 32'h00000000;
BRAM[2164]<= 32'h7E000000;
BRAM[2165]<= 32'h08081022;
BRAM[2166]<= 32'h00007E44;
BRAM[2167]<= 32'h00000000;
BRAM[2168]<= 32'h00000000;
BRAM[2169]<= 32'h00000000;
BRAM[2170]<= 32'hFF000000;
BRAM[2171]<= 32'h00000000;
BRAM[2172]<= 32'h18180000;
BRAM[2173]<= 32'h00000000;
BRAM[2174]<= 32'h00001818;
BRAM[2175]<= 32'h40000000;
BRAM[2176]<= 32'h04081020;
BRAM[2177]<= 32'h10080402;
BRAM[2178]<= 32'h00004020;
BRAM[2179]<= 32'h00000000;
BRAM[2180]<= 32'h00000000;
BRAM[2181]<= 32'h00000000;
BRAM[2182]<= 32'h00000000;
BRAM[2183]<= 32'h00000000;
BRAM[2184]<= 32'h10101000;
BRAM[2185]<= 32'h101010FE;
BRAM[2186]<= 32'h00000000;
BRAM[2187]<= 32'h00000000;
BRAM[2188]<= 32'h00000000;
BRAM[2189]<= 32'h0000007E;
BRAM[2190]<= 32'h00000000;
BRAM[2191]<= 32'h00000000;
BRAM[2192]<= 32'h00000000;
BRAM[2193]<= 32'h00000000;
BRAM[2194]<= 32'h00000000;
BRAM[2195]<= 32'h00000000;
BRAM[2196]<= 32'h00000000;
BRAM[2197]<= 32'h00000000;
BRAM[2198]<= 32'h00000000;
BRAM[2199]<= 32'h00000000;
BRAM[2200]<= 32'h00000000;
BRAM[2201]<= 32'h00003000;
BRAM[2202]<= 32'h00000000;
BRAM[2203]<= 32'h00000000;
BRAM[2204]<= 32'h00000000;
BRAM[2205]<= 32'h00000000;
BRAM[2206]<= 32'h00000000;
BRAM[2207]<= 32'h00000000;
BRAM[2208]<= 32'h00000000;
BRAM[2209]<= 32'h00000000;
BRAM[2210]<= 32'h00000000;
BRAM[2211]<= 32'h00003000;
BRAM[2212]<= 32'h003C0000;
BRAM[2213]<= 32'h00000000;
BRAM[2214]<= 32'h01000000;
BRAM[2215]<= 32'h000000C0;
BRAM[2216]<= 32'h00000006;
BRAM[2217]<= 32'h00000000;
BRAM[2218]<= 32'h01070000;
BRAM[2219]<= 32'h00F000E0;
BRAM[2220]<= 32'h00000000;
BRAM[2221]<= 32'h00003001;
BRAM[2222]<= 32'h00FE0000;
BRAM[2223]<= 32'h00000000;
BRAM[2224]<= 32'hC3011C00;
BRAM[2225]<= 32'h000000F0;
BRAM[2226]<= 32'h00000004;
BRAM[2227]<= 32'h00800C00;
BRAM[2228]<= 32'h070F0018;
BRAM[2229]<= 32'h00F803F8;
BRAM[2230]<= 32'h00000000;
BRAM[2231]<= 32'h03003001;
BRAM[2232]<= 32'h00FE0100;
BRAM[2233]<= 32'h00000000;
BRAM[2234]<= 32'hC7011C00;
BRAM[2235]<= 32'h000000F0;
BRAM[2236]<= 32'h4800000C;
BRAM[2237]<= 32'h03C00D00;
BRAM[2238]<= 32'h0F1F0018;
BRAM[2239]<= 32'h00F807F8;
BRAM[2240]<= 32'h60100000;
BRAM[2241]<= 32'h1F00B801;
BRAM[2242]<= 32'h00C60300;
BRAM[2243]<= 32'h00000000;
BRAM[2244]<= 32'hC7010C00;
BRAM[2245]<= 32'h80010078;
BRAM[2246]<= 32'hC800000C;
BRAM[2247]<= 32'h03800D00;
BRAM[2248]<= 32'h1E3B0018;
BRAM[2249]<= 32'h01100F3C;
BRAM[2250]<= 32'h60100007;
BRAM[2251]<= 32'h3F00F803;
BRAM[2252]<= 32'h00800300;
BRAM[2253]<= 32'h00000C00;
BRAM[2254]<= 32'hC2030E00;
BRAM[2255]<= 32'h80010038;
BRAM[2256]<= 32'hC800000D;
BRAM[2257]<= 32'h03800D00;
BRAM[2258]<= 32'h1C30001C;
BRAM[2259]<= 32'h01000E1E;
BRAM[2260]<= 32'h6038009F;
BRAM[2261]<= 32'hFC00F007;
BRAM[2262]<= 32'h00000700;
BRAM[2263]<= 32'h00000C00;
BRAM[2264]<= 32'hC0030E00;
BRAM[2265]<= 32'h80630018;
BRAM[2266]<= 32'h9B01800F;
BRAM[2267]<= 32'h03606F00;
BRAM[2268]<= 32'h38300008;
BRAM[2269]<= 32'h03001C0E;
BRAM[2270]<= 32'h6038009F;
BRAM[2271]<= 32'hFC00B007;
BRAM[2272]<= 32'h00000600;
BRAM[2273]<= 32'h00000C00;
BRAM[2274]<= 32'hC0030E00;
BRAM[2275]<= 32'h00730018;
BRAM[2276]<= 32'h9F01001F;
BRAM[2277]<= 32'h03E07F00;
BRAM[2278]<= 32'h38700000;
BRAM[2279]<= 32'h03001806;
BRAM[2280]<= 32'h601C0092;
BRAM[2281]<= 32'h1C003001;
BRAM[2282]<= 32'h00000E00;
BRAM[2283]<= 32'h00000C00;
BRAM[2284]<= 32'hC0030F00;
BRAM[2285]<= 32'h00730018;
BRAM[2286]<= 32'hDE011C1E;
BRAM[2287]<= 32'h03C06F00;
BRAM[2288]<= 32'h3070000E;
BRAM[2289]<= 32'h01003807;
BRAM[2290]<= 32'h60080096;
BRAM[2291]<= 32'h0C00F001;
BRAM[2292]<= 32'h1F000E00;
BRAM[2293]<= 32'h101FCC0C;
BRAM[2294]<= 32'hC0070F60;
BRAM[2295]<= 32'h00E60038;
BRAM[2296]<= 32'h7C037E16;
BRAM[2297]<= 32'h03806F00;
BRAM[2298]<= 32'h3070003F;
BRAM[2299]<= 32'h00003807;
BRAM[2300]<= 32'h60000096;
BRAM[2301]<= 32'h0C00B001;
BRAM[2302]<= 32'h3F000E00;
BRAM[2303]<= 32'h383FCF8D;
BRAM[2304]<= 32'hC0060B60;
BRAM[2305]<= 32'h00C60030;
BRAM[2306]<= 32'hF903FE07;
BRAM[2307]<= 32'h03806C00;
BRAM[2308]<= 32'h70308039;
BRAM[2309]<= 32'h00003007;
BRAM[2310]<= 32'h60000016;
BRAM[2311]<= 32'h0F003001;
BRAM[2312]<= 32'h7B000CC0;
BRAM[2313]<= 32'h9833FF8F;
BRAM[2314]<= 32'hC0060BE0;
BRAM[2315]<= 32'hE0C70070;
BRAM[2316]<= 32'hF907EE0F;
BRAM[2317]<= 32'h07C06D00;
BRAM[2318]<= 32'h703880F9;
BRAM[2319]<= 32'h00003007;
BRAM[2320]<= 32'h7C000036;
BRAM[2321]<= 32'h1F00F001;
BRAM[2322]<= 32'h61000CC0;
BRAM[2323]<= 32'h9C31FFCF;
BRAM[2324]<= 32'hC18E1BC0;
BRAM[2325]<= 32'hF08F01E0;
BRAM[2326]<= 32'hB907EE1F;
BRAM[2327]<= 32'h1F802D80;
BRAM[2328]<= 32'h703880FF;
BRAM[2329]<= 32'h00003007;
BRAM[2330]<= 32'hFC30003F;
BRAM[2331]<= 32'h7F00B001;
BRAM[2332]<= 32'hE1000CE0;
BRAM[2333]<= 32'h8C610CCE;
BRAM[2334]<= 32'hC38C19C0;
BRAM[2335]<= 32'hF0BE01C0;
BRAM[2336]<= 32'h0F0F6C7E;
BRAM[2337]<= 32'h1F802B80;
BRAM[2338]<= 32'h701C80FF;
BRAM[2339]<= 32'h01003003;
BRAM[2340]<= 32'hFCF38033;
BRAM[2341]<= 32'hFF013C01;
BRAM[2342]<= 32'hC0000CC0;
BRAM[2343]<= 32'h8D610CCE;
BRAM[2344]<= 32'hC38C1980;
BRAM[2345]<= 32'h60F801F0;
BRAM[2346]<= 32'hCF067CFF;
BRAM[2347]<= 32'h1F002A80;
BRAM[2348]<= 32'h701C00EC;
BRAM[2349]<= 32'h03003007;
BRAM[2350]<= 32'hE0F781B3;
BRAM[2351]<= 32'hCC07FE01;
BRAM[2352]<= 32'hC0000C00;
BRAM[2353]<= 32'h87610CCC;
BRAM[2354]<= 32'hC08C1980;
BRAM[2355]<= 32'h60980370;
BRAM[2356]<= 32'hE0057C6F;
BRAM[2357]<= 32'h1B002800;
BRAM[2358]<= 32'h700E00AE;
BRAM[2359]<= 32'h0F003007;
BRAM[2360]<= 32'hE0F7018E;
BRAM[2361]<= 32'h0C02F003;
BRAM[2362]<= 32'hC0000C00;
BRAM[2363]<= 32'h877F0CCC;
BRAM[2364]<= 32'hC0D8990F;
BRAM[2365]<= 32'h60980138;
BRAM[2366]<= 32'h6003780B;
BRAM[2367]<= 32'h07E00700;
BRAM[2368]<= 32'h700E0020;
BRAM[2369]<= 32'h1F003007;
BRAM[2370]<= 32'h60F0011F;
BRAM[2371]<= 32'h0C00F00F;
BRAM[2372]<= 32'hC0000E00;
BRAM[2373]<= 32'h877F0CCC;
BRAM[2374]<= 32'hC0D8980F;
BRAM[2375]<= 32'h60FF0118;
BRAM[2376]<= 32'hFB030019;
BRAM[2377]<= 32'h06E00F00;
BRAM[2378]<= 32'h70070060;
BRAM[2379]<= 32'h1F003807;
BRAM[2380]<= 32'h60200037;
BRAM[2381]<= 32'h0C00301F;
BRAM[2382]<= 32'hC0000E00;
BRAM[2383]<= 32'h076C0CCC;
BRAM[2384]<= 32'hC0D8180F;
BRAM[2385]<= 32'h60DB0118;
BRAM[2386]<= 32'hFB030018;
BRAM[2387]<= 32'h0E603F00;
BRAM[2388]<= 32'h7007000E;
BRAM[2389]<= 32'h13003806;
BRAM[2390]<= 32'h60240036;
BRAM[2391]<= 32'h0C00D802;
BRAM[2392]<= 32'hC0000E00;
BRAM[2393]<= 32'h0F600CCC;
BRAM[2394]<= 32'hC0F81800;
BRAM[2395]<= 32'h60DB0118;
BRAM[2396]<= 32'h5F03E039;
BRAM[2397]<= 32'h1E603F00;
BRAM[2398]<= 32'h3003003E;
BRAM[2399]<= 32'h03003806;
BRAM[2400]<= 32'h6024003E;
BRAM[2401]<= 32'h0C00DC06;
BRAM[2402]<= 32'hC0000700;
BRAM[2403]<= 32'h0D600CCC;
BRAM[2404]<= 32'hC0701880;
BRAM[2405]<= 32'h60990118;
BRAM[2406]<= 32'h7C03F027;
BRAM[2407]<= 32'h3E603F00;
BRAM[2408]<= 32'h3807007C;
BRAM[2409]<= 32'h03001C0E;
BRAM[2410]<= 32'h606C009E;
BRAM[2411]<= 32'h0C00FC06;
BRAM[2412]<= 32'hE0000700;
BRAM[2413]<= 32'h1D601CCC;
BRAM[2414]<= 32'hC0701880;
BRAM[2415]<= 32'h60980138;
BRAM[2416]<= 32'hFC037006;
BRAM[2417]<= 32'h7A403FC0;
BRAM[2418]<= 32'h3807007C;
BRAM[2419]<= 32'h03001C0C;
BRAM[2420]<= 32'h6068009E;
BRAM[2421]<= 32'h0C00F607;
BRAM[2422]<= 32'h61840300;
BRAM[2423]<= 32'h19701C8E;
BRAM[2424]<= 32'hE47018C0;
BRAM[2425]<= 32'h60F80138;
BRAM[2426]<= 32'h5803B006;
BRAM[2427]<= 32'h72E03FC0;
BRAM[2428]<= 32'h1C060018;
BRAM[2429]<= 32'h03100E1C;
BRAM[2430]<= 32'h6078008E;
BRAM[2431]<= 32'h0C00C70F;
BRAM[2432]<= 32'h73EE0300;
BRAM[2433]<= 32'h98390C8E;
BRAM[2434]<= 32'hE77038C0;
BRAM[2435]<= 32'h60F801F0;
BRAM[2436]<= 32'h5802B007;
BRAM[2437]<= 32'h22F83FC0;
BRAM[2438]<= 32'h1F7E001C;
BRAM[2439]<= 32'h03F80F78;
BRAM[2440]<= 32'h6078008F;
BRAM[2441]<= 32'h0C80C718;
BRAM[2442]<= 32'h7FFE0100;
BRAM[2443]<= 32'hB83F0E8E;
BRAM[2444]<= 32'hE72038E0;
BRAM[2445]<= 32'hE0FC00E0;
BRAM[2446]<= 32'h58023007;
BRAM[2447]<= 32'h06F83FC0;
BRAM[2448]<= 32'h0F7C801F;
BRAM[2449]<= 32'h03F807F8;
BRAM[2450]<= 32'h6030001F;
BRAM[2451]<= 32'h0CC0D338;
BRAM[2452]<= 32'h3FFC0000;
BRAM[2453]<= 32'h301F0E0E;
BRAM[2454]<= 32'hE7003860;
BRAM[2455]<= 32'hC0BE00E0;
BRAM[2456]<= 32'h58023006;
BRAM[2457]<= 32'h0EF87FC0;
BRAM[2458]<= 32'h077880FF;
BRAM[2459]<= 32'h03F003E0;
BRAM[2460]<= 32'h6030C079;
BRAM[2461]<= 32'h1C00F831;
BRAM[2462]<= 32'h0C380000;
BRAM[2463]<= 32'h000E0600;
BRAM[2464]<= 32'h03000000;
BRAM[2465]<= 32'hC0130080;
BRAM[2466]<= 32'hE8033006;
BRAM[2467]<= 32'h0F08F0C1;
BRAM[2468]<= 32'h013080F1;
BRAM[2469]<= 32'h02E00080;
BRAM[2470]<= 32'h6030F071;
BRAM[2471]<= 32'hF800F807;
BRAM[2472]<= 32'h00000000;
BRAM[2473]<= 32'h00000000;
BRAM[2474]<= 32'h00000000;
BRAM[2475]<= 32'hC0010000;
BRAM[2476]<= 32'hEF02B007;
BRAM[2477]<= 32'h0600C0C1;
BRAM[2478]<= 32'h00000080;
BRAM[2479]<= 32'h02000000;
BRAM[2480]<= 32'h6000F801;
BRAM[2481]<= 32'h78000007;
BRAM[2482]<= 32'h00000000;
BRAM[2483]<= 32'h00000000;
BRAM[2484]<= 32'h00000000;
BRAM[2485]<= 32'hC0000000;
BRAM[2486]<= 32'hEF00F007;
BRAM[2487]<= 32'h020000C0;
BRAM[2488]<= 32'h00000000;
BRAM[2489]<= 32'h00000000;
BRAM[2490]<= 32'h6000F800;
BRAM[2491]<= 32'h18000000;
BRAM[2492]<= 32'h00000000;
BRAM[2493]<= 32'h00000000;
BRAM[2494]<= 32'h00000000;
BRAM[2495]<= 32'h00000000;
BRAM[2496]<= 32'h60007002;
BRAM[2497]<= 32'h00000000;
BRAM[2498]<= 32'h00000000;
BRAM[2499]<= 32'h00000000;
BRAM[2500]<= 32'h60000000;
BRAM[2501]<= 32'h00000000;
BRAM[2502]<= 32'h00000000;
BRAM[2503]<= 32'h00000000;
BRAM[2504]<= 32'h00000000;
BRAM[2505]<= 32'h00000000;
BRAM[2506]<= 32'h00007000;
BRAM[2507]<= 32'h00000000;
BRAM[2508]<= 32'h00000000;
BRAM[2509]<= 32'h00000000;
BRAM[2510]<= 32'h60000000;
BRAM[2511]<= 32'hFFFFFFFF;
BRAM[2512]<= 32'hFFFFFFFF;
BRAM[2513]<= 32'hFFFFFFFF;
BRAM[2514]<= 32'hFFFFFFFF;
BRAM[2515]<= 32'hFFFFFFFF;
BRAM[2516]<= 32'hFFFFFFFF;
BRAM[2517]<= 32'hFFAA6AFF;
BRAM[2518]<= 32'hFFFFFFFF;
BRAM[2519]<= 32'hFFFFFFFF;
BRAM[2520]<= 32'hFFFFFFFF;
BRAM[2521]<= 32'hFFFFFFFF;
BRAM[2522]<= 32'hFFFFFFFF;
BRAM[2523]<= 32'hFFFFFFFF;
BRAM[2524]<= 32'hFFFFFFFF;
BRAM[2525]<= 32'hFFFFFFFF;
BRAM[2526]<= 32'hFFFFFFFF;
BRAM[2527]<= 32'hFFFFFFFF;
BRAM[2528]<= 32'hFFFFFFFF;
BRAM[2529]<= 32'hAAFAFFFF;
BRAM[2530]<= 32'hFFFFABAA;
BRAM[2531]<= 32'hFFFFFFFF;
BRAM[2532]<= 32'hFFFFFFFF;
BRAM[2533]<= 32'hFFFFFFFF;
BRAM[2534]<= 32'hFFFFFFFF;
BRAM[2535]<= 32'hFFFFFFFF;
BRAM[2536]<= 32'hFFFFFFFF;
BRAM[2537]<= 32'hFFFFFFFF;
BRAM[2538]<= 32'hFFFFFFFF;
BRAM[2539]<= 32'hFFFFFFFF;
BRAM[2540]<= 32'hFFFFFFFF;
BRAM[2541]<= 32'hFFFFFFFF;
BRAM[2542]<= 32'hAAAAAAAA;
BRAM[2543]<= 32'hFFFFFFBF;
BRAM[2544]<= 32'hFFFFFFFF;
BRAM[2545]<= 32'hFFFFFFFF;
BRAM[2546]<= 32'hFFFFFFFF;
BRAM[2547]<= 32'hFFFFFFFF;
BRAM[2548]<= 32'hFFFFFFFF;
BRAM[2549]<= 32'hFFFFFFFF;
BRAM[2550]<= 32'hFFFFFFFF;
BRAM[2551]<= 32'hFFFFFFFF;
BRAM[2552]<= 32'hFFFFFFFF;
BRAM[2553]<= 32'hFFFFFFFF;
BRAM[2554]<= 32'hAAAAFAFF;
BRAM[2555]<= 32'hFFAFAAAA;
BRAM[2556]<= 32'hFFFFFFFF;
BRAM[2557]<= 32'hFFFFFFFF;
BRAM[2558]<= 32'hFFFFFFFF;
BRAM[2559]<= 32'hFFFFFFFF;
BRAM[2560]<= 32'hFFFFFFFF;
BRAM[2561]<= 32'hFFFFFFFF;
BRAM[2562]<= 32'hFFFFFFFF;
BRAM[2563]<= 32'hFFFFFFFF;
BRAM[2564]<= 32'hFFFFFFFF;
BRAM[2565]<= 32'hFFFFFFFF;
BRAM[2566]<= 32'hAAFFFFFF;
BRAM[2567]<= 32'hAAAAAAAA;
BRAM[2568]<= 32'hFFFFFFAA;
BRAM[2569]<= 32'hFFFFFFFF;
BRAM[2570]<= 32'hFFFFFFFF;
BRAM[2571]<= 32'hFFFFFFFF;
BRAM[2572]<= 32'hFFFFFFFF;
BRAM[2573]<= 32'hFFFFFFFF;
BRAM[2574]<= 32'hFFFFFFFF;
BRAM[2575]<= 32'hFFFFFFFF;
BRAM[2576]<= 32'hFFFFFFFF;
BRAM[2577]<= 32'hFFFFFFFF;
BRAM[2578]<= 32'hFFFFFFFF;
BRAM[2579]<= 32'hAAAAAAFE;
BRAM[2580]<= 32'hAFAAAAAA;
BRAM[2581]<= 32'hFFFFFFFF;
BRAM[2582]<= 32'hFFFFFFFF;
BRAM[2583]<= 32'hFFFFFFFF;
BRAM[2584]<= 32'hFFFFFFFF;
BRAM[2585]<= 32'hFFFFFFFF;
BRAM[2586]<= 32'hFFFFFFFF;
BRAM[2587]<= 32'hFFFFFFFF;
BRAM[2588]<= 32'hFFFFFFFF;
BRAM[2589]<= 32'hFFFFFFFF;
BRAM[2590]<= 32'hFFFFFFFF;
BRAM[2591]<= 32'hAAEAFFFF;
BRAM[2592]<= 32'hAAAAAAAA;
BRAM[2593]<= 32'hFFFFAAAA;
BRAM[2594]<= 32'hFFFFFFFF;
BRAM[2595]<= 32'hFFFFFFFF;
BRAM[2596]<= 32'hFFFFFFFF;
BRAM[2597]<= 32'hFFFFFFFF;
BRAM[2598]<= 32'hFFFFFFFF;
BRAM[2599]<= 32'hFFFFFFFF;
BRAM[2600]<= 32'hFFFFFFFF;
BRAM[2601]<= 32'hFFFFFFFF;
BRAM[2602]<= 32'hFFFFFFFF;
BRAM[2603]<= 32'hFEFFFFFF;
BRAM[2604]<= 32'hAAAAAAAA;
BRAM[2605]<= 32'hAAAAAAAA;
BRAM[2606]<= 32'hFFFFFFBF;
BRAM[2607]<= 32'hFFFFFFFF;
BRAM[2608]<= 32'hFFFFFFFF;
BRAM[2609]<= 32'hFFFFFFFF;
BRAM[2610]<= 32'hFFFFFFFF;
BRAM[2611]<= 32'hFFFFFFFF;
BRAM[2612]<= 32'hFFFFFFFF;
BRAM[2613]<= 32'hFFFFFFFF;
BRAM[2614]<= 32'hFFFFFFFF;
BRAM[2615]<= 32'hFFFFFFFF;
BRAM[2616]<= 32'hAAAAEAFF;
BRAM[2617]<= 32'hAAAAAAAA;
BRAM[2618]<= 32'hFFABAAAA;
BRAM[2619]<= 32'hFFFFFFFF;
BRAM[2620]<= 32'hFFFFFFFF;
BRAM[2621]<= 32'hFFFFFFFF;
BRAM[2622]<= 32'hFFFFFFFF;
BRAM[2623]<= 32'hFFFFFFFF;
BRAM[2624]<= 32'hFFFFFFFF;
BRAM[2625]<= 32'hFFFFFFFF;
BRAM[2626]<= 32'hFFFFFFFF;
BRAM[2627]<= 32'hFFFFFFFF;
BRAM[2628]<= 32'hAAFEFFFF;
BRAM[2629]<= 32'hAAAAAAAA;
BRAM[2630]<= 32'hAAAAAAAA;
BRAM[2631]<= 32'hFFFFBFAA;
BRAM[2632]<= 32'hFFFFFFFF;
BRAM[2633]<= 32'hFFFFFFFF;
BRAM[2634]<= 32'hFFFFFFFF;
BRAM[2635]<= 32'hFFFFFFFF;
BRAM[2636]<= 32'hFFFFFFFF;
BRAM[2637]<= 32'hFFFFFFFF;
BRAM[2638]<= 32'hFFFFFFFF;
BRAM[2639]<= 32'hFFFFFFFF;
BRAM[2640]<= 32'hFFFFFFFF;
BRAM[2641]<= 32'hAAAAAAEA;
BRAM[2642]<= 32'hAAAAAAAA;
BRAM[2643]<= 32'hABAAAAAA;
BRAM[2644]<= 32'hFFFFFFFF;
BRAM[2645]<= 32'hFFFFFFFF;
BRAM[2646]<= 32'hFFFFFFFF;
BRAM[2647]<= 32'hFFFFFFFF;
BRAM[2648]<= 32'hFFFFFFFF;
BRAM[2649]<= 32'hFFFFFFFF;
BRAM[2650]<= 32'hFFFFFFFF;
BRAM[2651]<= 32'hFFFFFFFF;
BRAM[2652]<= 32'hFFFFFFFF;
BRAM[2653]<= 32'hAAAAFEFF;
BRAM[2654]<= 32'hAAAAAAAA;
BRAM[2655]<= 32'hAAAAAAAA;
BRAM[2656]<= 32'hFFBFAAAA;
BRAM[2657]<= 32'hFFFFFFFF;
BRAM[2658]<= 32'hFFFFFFFF;
BRAM[2659]<= 32'hFFFFFFFF;
BRAM[2660]<= 32'hFFFFFFFF;
BRAM[2661]<= 32'hFFFFFFFF;
BRAM[2662]<= 32'hFFFFFFFF;
BRAM[2663]<= 32'hFFFFFFFF;
BRAM[2664]<= 32'hFFFFFFFF;
BRAM[2665]<= 32'hEAFFFFFF;
BRAM[2666]<= 32'hAAAAAAAA;
BRAM[2667]<= 32'hAAAAAAAA;
BRAM[2668]<= 32'hAAAAAAAA;
BRAM[2669]<= 32'hFFFFFFAF;
BRAM[2670]<= 32'hFFFFFFFF;
BRAM[2671]<= 32'hFFFFFFFF;
BRAM[2672]<= 32'hFFFFFFFF;
BRAM[2673]<= 32'hFFFFFFFF;
BRAM[2674]<= 32'hFFFFFFFF;
BRAM[2675]<= 32'hFFFFFFFF;
BRAM[2676]<= 32'hFFFFFFFF;
BRAM[2677]<= 32'hFFFFFFFF;
BRAM[2678]<= 32'hAAAAEAFF;
BRAM[2679]<= 32'hAAAAAAAA;
BRAM[2680]<= 32'hAAAAAAAA;
BRAM[2681]<= 32'hFFAAAAAA;
BRAM[2682]<= 32'hFFFFFFFF;
BRAM[2683]<= 32'hFFFFFFFF;
BRAM[2684]<= 32'hFFFFFFFF;
BRAM[2685]<= 32'hFFFFFFFF;
BRAM[2686]<= 32'hFFFFFFFF;
BRAM[2687]<= 32'hFFFFFFFF;
BRAM[2688]<= 32'hFFFFFFFF;
BRAM[2689]<= 32'hFFFFFFFF;
BRAM[2690]<= 32'hFEFFFFFF;
BRAM[2691]<= 32'hAAAAAAAA;
BRAM[2692]<= 32'hAAAAAAAA;
BRAM[2693]<= 32'hAAAAAAAA;
BRAM[2694]<= 32'hFFFFAFAA;
BRAM[2695]<= 32'hFFFFFFFF;
BRAM[2696]<= 32'hFFFFFFFF;
BRAM[2697]<= 32'hFFFFFFFF;
BRAM[2698]<= 32'hFFFFFFFF;
BRAM[2699]<= 32'hFFFFFFFF;
BRAM[2700]<= 32'hFFFFFFFF;
BRAM[2701]<= 32'hFFFFFFFF;
BRAM[2702]<= 32'hFFFFFFFF;
BRAM[2703]<= 32'hAAEAFFFF;
BRAM[2704]<= 32'hAAAAAAAA;
BRAM[2705]<= 32'hAAAAAAAA;
BRAM[2706]<= 32'hAAAAAAAA;
BRAM[2707]<= 32'hFFFFFFFF;
BRAM[2708]<= 32'hFFFFFFFF;
BRAM[2709]<= 32'hFFFFFFFF;
BRAM[2710]<= 32'hFFFFFFFF;
BRAM[2711]<= 32'hFFFFFFFF;
BRAM[2712]<= 32'hFFFFFFFF;
BRAM[2713]<= 32'hFFFFFFFF;
BRAM[2714]<= 32'hFFFFFFFF;
BRAM[2715]<= 32'hFFAFFAFF;
BRAM[2716]<= 32'hAAAAAAFE;
BRAM[2717]<= 32'hAAAAAAAA;
BRAM[2718]<= 32'hAAAAAAAA;
BRAM[2719]<= 32'hFFBFAAAA;
BRAM[2720]<= 32'hFFFFFFFF;
BRAM[2721]<= 32'hFFFFFFFF;
BRAM[2722]<= 32'hFFFFFFFF;
BRAM[2723]<= 32'hFFFFFFFF;
BRAM[2724]<= 32'hFFFFFFFF;
BRAM[2725]<= 32'hFFFFFFFF;
BRAM[2726]<= 32'hFFFFFFFF;
BRAM[2727]<= 32'hAAFFFFFF;
BRAM[2728]<= 32'hAAFFFFAA;
BRAM[2729]<= 32'hAAAAAAAA;
BRAM[2730]<= 32'hAAAAAAAA;
BRAM[2731]<= 32'hAAAAAAAA;
BRAM[2732]<= 32'hFFFFFFAB;
BRAM[2733]<= 32'hFFFFFFFF;
BRAM[2734]<= 32'hFFFFFFFF;
BRAM[2735]<= 32'hFFFFFFFF;
BRAM[2736]<= 32'hFFFFFFFF;
BRAM[2737]<= 32'hFFFFFFFF;
BRAM[2738]<= 32'hFFFFFFFF;
BRAM[2739]<= 32'hFFFFFFFF;
BRAM[2740]<= 32'hAFAAAAFE;
BRAM[2741]<= 32'hAAAAFAFF;
BRAM[2742]<= 32'hAAAAAAAA;
BRAM[2743]<= 32'hAAAAAAAA;
BRAM[2744]<= 32'hBFAAAAAA;
BRAM[2745]<= 32'hFFFFFFFF;
BRAM[2746]<= 32'hFFFFFFFF;
BRAM[2747]<= 32'hFFFFFFFF;
BRAM[2748]<= 32'hFFFFFFFF;
BRAM[2749]<= 32'hFFFFFFFF;
BRAM[2750]<= 32'hFFFFFFFF;
BRAM[2751]<= 32'hFFFFFFFF;
BRAM[2752]<= 32'hAAEAFFFF;
BRAM[2753]<= 32'hFFFFAAAA;
BRAM[2754]<= 32'hAAAAAAAA;
BRAM[2755]<= 32'hAAAAAAAA;
BRAM[2756]<= 32'hAAAAAAAA;
BRAM[2757]<= 32'hFFFFABAA;
BRAM[2758]<= 32'hFFFFFFFF;
BRAM[2759]<= 32'hFFFFFFFF;
BRAM[2760]<= 32'hFFFFFFFF;
BRAM[2761]<= 32'hFFFFFFFF;
BRAM[2762]<= 32'hFFFFFFFF;
BRAM[2763]<= 32'hFFFFFFFF;
BRAM[2764]<= 32'hFEFFFFFF;
BRAM[2765]<= 32'hAAAAAAAA;
BRAM[2766]<= 32'hAAFAFFAF;
BRAM[2767]<= 32'hAAAAAAAA;
BRAM[2768]<= 32'hAAAAAAAA;
BRAM[2769]<= 32'hAAAAAAAA;
BRAM[2770]<= 32'hFFFFFFBF;
BRAM[2771]<= 32'hFFFFFFFF;
BRAM[2772]<= 32'hFFFFFFFF;
BRAM[2773]<= 32'hFFFFFFFF;
BRAM[2774]<= 32'hFFFFFFFF;
BRAM[2775]<= 32'hFFFFFFFF;
BRAM[2776]<= 32'hFFFFFFFF;
BRAM[2777]<= 32'hAAAAEAFF;
BRAM[2778]<= 32'hFFABAAAA;
BRAM[2779]<= 32'hAAAAAAFF;
BRAM[2780]<= 32'hAAAAAAAA;
BRAM[2781]<= 32'hAAAAAAAA;
BRAM[2782]<= 32'hFFAFAAAA;
BRAM[2783]<= 32'hFFFFFFFF;
BRAM[2784]<= 32'hFFFFFFFF;
BRAM[2785]<= 32'hFFFFFFFF;
BRAM[2786]<= 32'hFFFFFFFF;
BRAM[2787]<= 32'hFFFFFFFF;
BRAM[2788]<= 32'hFFFFFFFF;
BRAM[2789]<= 32'hAAFEFFFF;
BRAM[2790]<= 32'hAAAAAAAA;
BRAM[2791]<= 32'hEAFFBFAA;
BRAM[2792]<= 32'hAAAAAAAA;
BRAM[2793]<= 32'hAAAAAAAA;
BRAM[2794]<= 32'hAAAAAAAA;
BRAM[2795]<= 32'hFFFFFFAA;
BRAM[2796]<= 32'hFFFFFFFF;
BRAM[2797]<= 32'hFFFFFFFF;
BRAM[2798]<= 32'hFFFFFFFF;
BRAM[2799]<= 32'hFFFFFFFF;
BRAM[2800]<= 32'hFFFFFFFF;
BRAM[2801]<= 32'hFFFFFFFF;
BRAM[2802]<= 32'hAAAAAAEA;
BRAM[2803]<= 32'hABAAAAAA;
BRAM[2804]<= 32'hAAAAFEFF;
BRAM[2805]<= 32'hAAAAAAAA;
BRAM[2806]<= 32'hAAAAAAAA;
BRAM[2807]<= 32'hAFAAAAAA;
BRAM[2808]<= 32'hFFFFFFFF;
BRAM[2809]<= 32'hFFFFFFFF;
BRAM[2810]<= 32'hFFFFFFFF;
BRAM[2811]<= 32'hFFFFFFFF;
BRAM[2812]<= 32'hFFFFFFFF;
BRAM[2813]<= 32'hFFFFFFFF;
BRAM[2814]<= 32'hAAAAFFFF;
BRAM[2815]<= 32'hAAAAAAAA;
BRAM[2816]<= 32'hFFBFAAAA;
BRAM[2817]<= 32'hAAAAAAEA;
BRAM[2818]<= 32'hAAAAAAAA;
BRAM[2819]<= 32'hAAAAAAAA;
BRAM[2820]<= 32'hFFFFAAAA;
BRAM[2821]<= 32'hFFFFFFFF;
BRAM[2822]<= 32'hFFFFFFFF;
BRAM[2823]<= 32'hFFFFFFFF;
BRAM[2824]<= 32'hFFFFFFFF;
BRAM[2825]<= 32'hFFFFFFFF;
BRAM[2826]<= 32'hFAFFFFFF;
BRAM[2827]<= 32'hAAAAAAAA;
BRAM[2828]<= 32'hAAAAAAAA;
BRAM[2829]<= 32'hAAFEFFAF;
BRAM[2830]<= 32'hAAAAAAAA;
BRAM[2831]<= 32'hAAAAAAAA;
BRAM[2832]<= 32'hAAAAAAAA;
BRAM[2833]<= 32'hFFFFFFBF;
BRAM[2834]<= 32'hFFFFFFFF;
BRAM[2835]<= 32'hFFFFFFFF;
BRAM[2836]<= 32'hFFFFFFFF;
BRAM[2837]<= 32'hFFFFFFFF;
BRAM[2838]<= 32'hFFFFFFFF;
BRAM[2839]<= 32'hAAAAAAFF;
BRAM[2840]<= 32'hAAAAAAAA;
BRAM[2841]<= 32'hFFAAAAAA;
BRAM[2842]<= 32'hAAAAAAFF;
BRAM[2843]<= 32'hAAAAAAAA;
BRAM[2844]<= 32'hAAAAAAAA;
BRAM[2845]<= 32'hFFABAAAA;
BRAM[2846]<= 32'hFFFFFFFF;
BRAM[2847]<= 32'hFFFFFFFF;
BRAM[2848]<= 32'hFFFFFFFF;
BRAM[2849]<= 32'hFFFFFFFF;
BRAM[2850]<= 32'hFFFFFFFF;
BRAM[2851]<= 32'hAAFAFFFF;
BRAM[2852]<= 32'hAAAAAAAA;
BRAM[2853]<= 32'hAAAAAAAA;
BRAM[2854]<= 32'hFFFFAFAA;
BRAM[2855]<= 32'hAAAAAAFE;
BRAM[2856]<= 32'hAAAAAAAA;
BRAM[2857]<= 32'hAAAAAAAA;
BRAM[2858]<= 32'hFFFFBFAA;
BRAM[2859]<= 32'hFFFFFFFF;
BRAM[2860]<= 32'hFFFFFFFF;
BRAM[2861]<= 32'hFFFFFFFF;
BRAM[2862]<= 32'hFFFFFFFF;
BRAM[2863]<= 32'hFFFFFFFF;
BRAM[2864]<= 32'hAAAAAAAA;
BRAM[2865]<= 32'hAAAAAAAA;
BRAM[2866]<= 32'hAAAAAAAA;
BRAM[2867]<= 32'hAAFFFFFF;
BRAM[2868]<= 32'hAAAAAAAA;
BRAM[2869]<= 32'hAAAAAAAA;
BRAM[2870]<= 32'hABAAAAAA;
BRAM[2871]<= 32'hFFFFFFFF;
BRAM[2872]<= 32'hFFFFFFFF;
BRAM[2873]<= 32'hFFFFFFFF;
BRAM[2874]<= 32'hFFFFFFFF;
BRAM[2875]<= 32'hFFFFFFFF;
BRAM[2876]<= 32'hAAAAFAFF;
BRAM[2877]<= 32'hAAAAAAAA;
BRAM[2878]<= 32'hAAAAAAAA;
BRAM[2879]<= 32'hFFFFAAAA;
BRAM[2880]<= 32'hAAAAEAFF;
BRAM[2881]<= 32'hAAAAAAAA;
BRAM[2882]<= 32'hAAAAAAAA;
BRAM[2883]<= 32'hFFBFAAAA;
BRAM[2884]<= 32'hFFFFFFFF;
BRAM[2885]<= 32'hFFFFFFFF;
BRAM[2886]<= 32'hFFFFFFFF;
BRAM[2887]<= 32'hFFFFFFFF;
BRAM[2888]<= 32'hEAFFFFFF;
BRAM[2889]<= 32'hAAAAAAAA;
BRAM[2890]<= 32'hAAAAAAAA;
BRAM[2891]<= 32'hAAAAAAAA;
BRAM[2892]<= 32'hEAFFFFFF;
BRAM[2893]<= 32'hAAAAAAAA;
BRAM[2894]<= 32'hAAAAAAAA;
BRAM[2895]<= 32'hAAAAAAAA;
BRAM[2896]<= 32'hFFFFFFAF;
BRAM[2897]<= 32'hFFFFFFFF;
BRAM[2898]<= 32'hFFFFFFFF;
BRAM[2899]<= 32'hFFFFFFFF;
BRAM[2900]<= 32'hFFFFFFFF;
BRAM[2901]<= 32'hAAAAAAFE;
BRAM[2902]<= 32'hAAAAAAAA;
BRAM[2903]<= 32'hAAAAAAAA;
BRAM[2904]<= 32'hFFBFAAAA;
BRAM[2905]<= 32'hAAAAEAFF;
BRAM[2906]<= 32'hAAAAAAAA;
BRAM[2907]<= 32'hAAAAAAAA;
BRAM[2908]<= 32'hFFAAAAAA;
BRAM[2909]<= 32'hFFFFFFFF;
BRAM[2910]<= 32'hFFFFFFFF;
BRAM[2911]<= 32'hFFFFFFFF;
BRAM[2912]<= 32'hFFFFFFFF;
BRAM[2913]<= 32'hAAEAFFFF;
BRAM[2914]<= 32'hAAAAAAAA;
BRAM[2915]<= 32'hAAAAAAAA;
BRAM[2916]<= 32'hAAAAAAAA;
BRAM[2917]<= 32'hFEFFFFFF;
BRAM[2918]<= 32'hAAAAAAAA;
BRAM[2919]<= 32'hAAAAAAAA;
BRAM[2920]<= 32'hAAAAAAAA;
BRAM[2921]<= 32'hFFFFAFAA;
BRAM[2922]<= 32'hFFFFFFFF;
BRAM[2923]<= 32'hFFFFFFFF;
BRAM[2924]<= 32'hFFFFFFFF;
BRAM[2925]<= 32'hFEFFFFFF;
BRAM[2926]<= 32'hAAAAAAAA;
BRAM[2927]<= 32'hAAAAAAAA;
BRAM[2928]<= 32'hAAAAAAAA;
BRAM[2929]<= 32'hFFFFAFAA;
BRAM[2930]<= 32'hAAEAFFFF;
BRAM[2931]<= 32'hAAAAAAAA;
BRAM[2932]<= 32'hAAAAAAAA;
BRAM[2933]<= 32'hABAAAAAA;
BRAM[2934]<= 32'hFFFFFFFF;
BRAM[2935]<= 32'hFFFFFFFF;
BRAM[2936]<= 32'hFFFFFFFF;
BRAM[2937]<= 32'hFFFFFFFF;
BRAM[2938]<= 32'hAAAAEAFF;
BRAM[2939]<= 32'hAAAAAAAA;
BRAM[2940]<= 32'hAAAAAAAA;
BRAM[2941]<= 32'hFFAAAAAA;
BRAM[2942]<= 32'hFFABAAFF;
BRAM[2943]<= 32'hAAAAAAFE;
BRAM[2944]<= 32'hAAAAAAAA;
BRAM[2945]<= 32'hAAAAAAAA;
BRAM[2946]<= 32'hFFFFABAA;
BRAM[2947]<= 32'hFFFFFFFF;
BRAM[2948]<= 32'hFFFFFFFF;
BRAM[2949]<= 32'hFFFFFFFF;
BRAM[2950]<= 32'hAAFEFFFF;
BRAM[2951]<= 32'hAAAAAAAA;
BRAM[2952]<= 32'hAAAAAAAA;
BRAM[2953]<= 32'hAAAAAAAA;
BRAM[2954]<= 32'hAAFAFFAF;
BRAM[2955]<= 32'hAAFFFFAA;
BRAM[2956]<= 32'hAAAAAAAA;
BRAM[2957]<= 32'hAAAAAAAA;
BRAM[2958]<= 32'hBFAAAAAA;
BRAM[2959]<= 32'hFFFFFFFF;
BRAM[2960]<= 32'hFFFFFFFF;
BRAM[2961]<= 32'hFFFFFFFF;
BRAM[2962]<= 32'hFFFFFFFF;
BRAM[2963]<= 32'hAAAAAAFA;
BRAM[2964]<= 32'hAAAAAAAA;
BRAM[2965]<= 32'hAAAAAAAA;
BRAM[2966]<= 32'hFFFFAAAA;
BRAM[2967]<= 32'hAFAAAAAA;
BRAM[2968]<= 32'hAAAAFAFF;
BRAM[2969]<= 32'hAAAAAAAA;
BRAM[2970]<= 32'hAAAAAAAA;
BRAM[2971]<= 32'hBFFEFFAB;
BRAM[2972]<= 32'hFFFFFFFF;
BRAM[2973]<= 32'hFFFFFFFF;
BRAM[2974]<= 32'hFFFFFFFF;
BRAM[2975]<= 32'hAAAAFFFF;
BRAM[2976]<= 32'hAAAAAAAA;
BRAM[2977]<= 32'hAAAAAAAA;
BRAM[2978]<= 32'hAFAAAAAA;
BRAM[2979]<= 32'hAAAAFEFF;
BRAM[2980]<= 32'hFFFFAAAA;
BRAM[2981]<= 32'hAAAAAAAA;
BRAM[2982]<= 32'hAAAAAAAA;
BRAM[2983]<= 32'hFFBFAAAA;
BRAM[2984]<= 32'hFFFFABEA;
BRAM[2985]<= 32'hFFFFFFFF;
BRAM[2986]<= 32'hFFFFFFFF;
BRAM[2987]<= 32'hFAFFFFFF;
BRAM[2988]<= 32'hAAAAAAAA;
BRAM[2989]<= 32'hAAAAAAAA;
BRAM[2990]<= 32'hAAAAAAAA;
BRAM[2991]<= 32'hEAFFFFAA;
BRAM[2992]<= 32'hAAAAAAAA;
BRAM[2993]<= 32'hAAFAFFAF;
BRAM[2994]<= 32'hAAAAAAAA;
BRAM[2995]<= 32'hABAAAAAA;
BRAM[2996]<= 32'hAAAAFEFF;
BRAM[2997]<= 32'hFFFFFFBF;
BRAM[2998]<= 32'hFFFFFFFF;
BRAM[2999]<= 32'hFFFFFFFF;
BRAM[3000]<= 32'hAAAAAAFF;
BRAM[3001]<= 32'hAAAAAAAA;
BRAM[3002]<= 32'hAAAAAAAA;
BRAM[3003]<= 32'hFFABAAAA;
BRAM[3004]<= 32'hAAAAAAFE;
BRAM[3005]<= 32'hFFABAAAA;
BRAM[3006]<= 32'hAAAAAAFF;
BRAM[3007]<= 32'hAAAAAAAA;
BRAM[3008]<= 32'hFAFFBFAA;
BRAM[3009]<= 32'hFFAFAAAA;
BRAM[3010]<= 32'hFFFFFFFF;
BRAM[3011]<= 32'hFFFFFFFF;
BRAM[3012]<= 32'hAAFAFFFF;
BRAM[3013]<= 32'hAAAAAAAA;
BRAM[3014]<= 32'hAAAAAAAA;
BRAM[3015]<= 32'hAAAAAAAA;
BRAM[3016]<= 32'hAAEAFFBF;
BRAM[3017]<= 32'hAAAAAAAA;
BRAM[3018]<= 32'hEAFFBFAA;
BRAM[3019]<= 32'hAAAAAAAA;
BRAM[3020]<= 32'hFFAAAAAA;
BRAM[3021]<= 32'hAAAAAAFF;
BRAM[3022]<= 32'hFFFFFFAA;
BRAM[3023]<= 32'hFFFFFFFF;
BRAM[3024]<= 32'hFFFFFFFF;
BRAM[3025]<= 32'hAAAAAAAA;
BRAM[3026]<= 32'hAAAAAAAA;
BRAM[3027]<= 32'hAAAAAAAA;
BRAM[3028]<= 32'hFEFFABAA;
BRAM[3029]<= 32'hAAAAAAAA;
BRAM[3030]<= 32'hABAAAAAA;
BRAM[3031]<= 32'hAAAAFEFF;
BRAM[3032]<= 32'hAAAAAAAA;
BRAM[3033]<= 32'hAAFAFFAF;
BRAM[3034]<= 32'hAFAAAAAA;
BRAM[3035]<= 32'hFFFFFFFF;
BRAM[3036]<= 32'hFFFFFFFF;
BRAM[3037]<= 32'hAAAAFAFF;
BRAM[3038]<= 32'hAAAAAAAA;
BRAM[3039]<= 32'hAAAAAAAA;
BRAM[3040]<= 32'hBFAAAAAA;
BRAM[3041]<= 32'hAAAAEAFF;
BRAM[3042]<= 32'hAAAAAAAA;
BRAM[3043]<= 32'hFFBFAAAA;
BRAM[3044]<= 32'hAAAAAAEA;
BRAM[3045]<= 32'hFFFFAAAA;
BRAM[3046]<= 32'hAAAAAAAA;
BRAM[3047]<= 32'hFFFFAAAA;
BRAM[3048]<= 32'hFFFFFFFF;
BRAM[3049]<= 32'hAAFFFFFF;
BRAM[3050]<= 32'hAAAAAAAA;
BRAM[3051]<= 32'hAAAAAAAA;
BRAM[3052]<= 32'hAAAAAAAA;
BRAM[3053]<= 32'hAAFEFFAB;
BRAM[3054]<= 32'hAAAAAAAA;
BRAM[3055]<= 32'hAAAAAAAA;
BRAM[3056]<= 32'hAAFEFFAB;
BRAM[3057]<= 32'hAFAAAAAA;
BRAM[3058]<= 32'hAAAAFAFF;
BRAM[3059]<= 32'hAAAAAAAA;
BRAM[3060]<= 32'hFFFFFFAF;
BRAM[3061]<= 32'hFFFFFFFF;
BRAM[3062]<= 32'hAAAAAAFE;
BRAM[3063]<= 32'hAAAAAAAA;
BRAM[3064]<= 32'hAAAAAAAA;
BRAM[3065]<= 32'hFFBFAAAA;
BRAM[3066]<= 32'hAAAAAAFA;
BRAM[3067]<= 32'hAAAAAAAA;
BRAM[3068]<= 32'hFFAAAAAA;
BRAM[3069]<= 32'hAAAAAAFF;
BRAM[3070]<= 32'hAAFFFFAA;
BRAM[3071]<= 32'hAAAAAAAA;
BRAM[3072]<= 32'hFFABAAAA;
BRAM[3073]<= 32'hFFFFFFFF;
BRAM[3074]<= 32'hAAEAFFFF;
BRAM[3075]<= 32'hAAAAAAAA;
BRAM[3076]<= 32'hAAAAAAAA;
BRAM[3077]<= 32'hABAAAAAA;
BRAM[3078]<= 32'hAAAAFFFF;
BRAM[3079]<= 32'hAAAAAAAA;
BRAM[3080]<= 32'hAAAAAAAA;
BRAM[3081]<= 32'hFAFFAFAA;
BRAM[3082]<= 32'hFFAFAAAA;
BRAM[3083]<= 32'hAAAAAAFA;
BRAM[3084]<= 32'hAAAAAAAA;
BRAM[3085]<= 32'hFFFFBFAA;
BRAM[3086]<= 32'hFEFFFFFF;
BRAM[3087]<= 32'hAAAAAAAA;
BRAM[3088]<= 32'hAAAAAAAA;
BRAM[3089]<= 32'hAAAAAAAA;
BRAM[3090]<= 32'hFAFFAFAA;
BRAM[3091]<= 32'hAAAAAAAA;
BRAM[3092]<= 32'hAAAAAAAA;
BRAM[3093]<= 32'hAAAAAAAA;
BRAM[3094]<= 32'hAAAAFFFF;
BRAM[3095]<= 32'hAAEAFFFF;
BRAM[3096]<= 32'hAAAAAAAA;
BRAM[3097]<= 32'hABAAAAAA;
BRAM[3098]<= 32'hFFFFFFFF;
BRAM[3099]<= 32'hAAAAEAFF;
BRAM[3100]<= 32'hAAAAAAAA;
BRAM[3101]<= 32'hAAAAAAAA;
BRAM[3102]<= 32'hFFFFAAAA;
BRAM[3103]<= 32'hAAAAAAFF;
BRAM[3104]<= 32'hAAAAAAAA;
BRAM[3105]<= 32'hAAAAAAAA;
BRAM[3106]<= 32'hFFAFAAAA;
BRAM[3107]<= 32'hFEFFFFFB;
BRAM[3108]<= 32'hAAAAAAAA;
BRAM[3109]<= 32'hAAAAAAAA;
BRAM[3110]<= 32'hFFBFAAAA;
BRAM[3111]<= 32'hAAFEFFFF;
BRAM[3112]<= 32'hAAAAAAAA;
BRAM[3113]<= 32'hAAAAAAAA;
BRAM[3114]<= 32'hBFAAAAAA;
BRAM[3115]<= 32'hAAFAFFFF;
BRAM[3116]<= 32'hAAAAAAAA;
BRAM[3117]<= 32'hAAAAAAAA;
BRAM[3118]<= 32'hAAAAAAAA;
BRAM[3119]<= 32'hFFFFFFAA;
BRAM[3120]<= 32'hAAAAEAFF;
BRAM[3121]<= 32'hAAAAAAAA;
BRAM[3122]<= 32'hAAAAAAAA;
BRAM[3123]<= 32'hFFFFFFAF;
BRAM[3124]<= 32'hAAAAAAFA;
BRAM[3125]<= 32'hAAAAAAAA;
BRAM[3126]<= 32'hAAAAAAAA;
BRAM[3127]<= 32'hFFFFFFAA;
BRAM[3128]<= 32'hAAAAAAAA;
BRAM[3129]<= 32'hAAAAAAAA;
BRAM[3130]<= 32'hAAAAAAAA;
BRAM[3131]<= 32'hBFAAAAAA;
BRAM[3132]<= 32'hAAFEFFFF;
BRAM[3133]<= 32'hAAAAAAAA;
BRAM[3134]<= 32'hAAAAAAAA;
BRAM[3135]<= 32'hFFAAAAAA;
BRAM[3136]<= 32'hAAEAFFFF;
BRAM[3137]<= 32'hAAAAAAAA;
BRAM[3138]<= 32'hAAAAAAAA;
BRAM[3139]<= 32'hFFABAAAA;
BRAM[3140]<= 32'hAAAAFFFF;
BRAM[3141]<= 32'hAAAAAAAA;
BRAM[3142]<= 32'hAAAAAAAA;
BRAM[3143]<= 32'hAAAAAAAA;
BRAM[3144]<= 32'hFFFFAFAA;
BRAM[3145]<= 32'hAAAAAAFE;
BRAM[3146]<= 32'hAAAAAAAA;
BRAM[3147]<= 32'hAAAAAAAA;
BRAM[3148]<= 32'hFFFFFFAA;
BRAM[3149]<= 32'hAAAAAAEA;
BRAM[3150]<= 32'hAAAAAAAA;
BRAM[3151]<= 32'hAAAAAAAA;
BRAM[3152]<= 32'hFFFFFFAB;
BRAM[3153]<= 32'hAAAAAAAA;
BRAM[3154]<= 32'hAAAAAAAA;
BRAM[3155]<= 32'hAAAAAAAA;
BRAM[3156]<= 32'hABAAAAAA;
BRAM[3157]<= 32'hAAFEFFFF;
BRAM[3158]<= 32'hAAAAAAAA;
BRAM[3159]<= 32'hAAAAAAAA;
BRAM[3160]<= 32'hBFAAAAAA;
BRAM[3161]<= 32'hAAEAFFFF;
BRAM[3162]<= 32'hAAAAAAAA;
BRAM[3163]<= 32'hAAAAAAAA;
BRAM[3164]<= 32'hFFABAAAA;
BRAM[3165]<= 32'hAAFAFFFF;
BRAM[3166]<= 32'hAAAAAAAA;
BRAM[3167]<= 32'hAAAAAAAA;
BRAM[3168]<= 32'hAAAAAAAA;
BRAM[3169]<= 32'hFFFFBFAA;
BRAM[3170]<= 32'hAAAAAAFA;
BRAM[3171]<= 32'hAAAAAAAA;
BRAM[3172]<= 32'hAAAAAAAA;
BRAM[3173]<= 32'hFFFFBFAA;
BRAM[3174]<= 32'hAAAAAAEA;
BRAM[3175]<= 32'hAAAAAAAA;
BRAM[3176]<= 32'hAAAAAAAA;
BRAM[3177]<= 32'hFFFFFFBF;
BRAM[3178]<= 32'hAAAAAAFF;
BRAM[3179]<= 32'hAAAAAAAA;
BRAM[3180]<= 32'hAAAAAAAA;
BRAM[3181]<= 32'hFFABAAAA;
BRAM[3182]<= 32'hAAEAFFFF;
BRAM[3183]<= 32'hAAAAAAAA;
BRAM[3184]<= 32'hAAAAAAAA;
BRAM[3185]<= 32'hFFAAAAAA;
BRAM[3186]<= 32'hAAEAFFFF;
BRAM[3187]<= 32'hAAAAAAAA;
BRAM[3188]<= 32'hAAAAAAAA;
BRAM[3189]<= 32'hFEFFABAA;
BRAM[3190]<= 32'hEAFFBFAA;
BRAM[3191]<= 32'hAAAAAAAA;
BRAM[3192]<= 32'hAAAAAAAA;
BRAM[3193]<= 32'hAAAAAAAA;
BRAM[3194]<= 32'hAAFAFFAF;
BRAM[3195]<= 32'hAAAAAAAA;
BRAM[3196]<= 32'hAAAAAAAA;
BRAM[3197]<= 32'hAAAAAAAA;
BRAM[3198]<= 32'hFFFFFFAB;
BRAM[3199]<= 32'hAAAAAAEA;
BRAM[3200]<= 32'hAAAAAAAA;
BRAM[3201]<= 32'hBFAAAAAA;
BRAM[3202]<= 32'hABAAEAFF;
BRAM[3203]<= 32'hAAAAFEFF;
BRAM[3204]<= 32'hAAAAAAAA;
BRAM[3205]<= 32'hAAAAAAAA;
BRAM[3206]<= 32'hFFFFAAAA;
BRAM[3207]<= 32'hAAAAAAAA;
BRAM[3208]<= 32'hAAAAAAAA;
BRAM[3209]<= 32'hAAAAAAAA;
BRAM[3210]<= 32'hFFBFAAAA;
BRAM[3211]<= 32'hBAEAFFFF;
BRAM[3212]<= 32'hAAAAAAAA;
BRAM[3213]<= 32'hAAAAAAAA;
BRAM[3214]<= 32'hAAFEFFAB;
BRAM[3215]<= 32'hFFBFAAAA;
BRAM[3216]<= 32'hAAAAAAEA;
BRAM[3217]<= 32'hAAAAAAAA;
BRAM[3218]<= 32'hAFAAAAAA;
BRAM[3219]<= 32'hAAAAFAFF;
BRAM[3220]<= 32'hAAAAAAAA;
BRAM[3221]<= 32'hAAAAAAAA;
BRAM[3222]<= 32'hABAAAAAA;
BRAM[3223]<= 32'hFFFFFFFF;
BRAM[3224]<= 32'hAAAABFEA;
BRAM[3225]<= 32'hAAAAAAAA;
BRAM[3226]<= 32'hFFBFAAAA;
BRAM[3227]<= 32'hAAAAAAEA;
BRAM[3228]<= 32'hAAFEFFAB;
BRAM[3229]<= 32'hAAAAAAAA;
BRAM[3230]<= 32'hAAAAAAAA;
BRAM[3231]<= 32'hAAFFFFAA;
BRAM[3232]<= 32'hAAAAAAAA;
BRAM[3233]<= 32'hAAAAAAAA;
BRAM[3234]<= 32'hAAAAAAAA;
BRAM[3235]<= 32'hFFFFAFAA;
BRAM[3236]<= 32'hBFEAFFFF;
BRAM[3237]<= 32'hAAAAAAFA;
BRAM[3238]<= 32'hABAAAAAA;
BRAM[3239]<= 32'hAAAAFFFF;
BRAM[3240]<= 32'hFFAAAAAA;
BRAM[3241]<= 32'hAAAAAAFF;
BRAM[3242]<= 32'hAAAAAAAA;
BRAM[3243]<= 32'hFFAFAAAA;
BRAM[3244]<= 32'hAAAAAAFA;
BRAM[3245]<= 32'hAAAAAAAA;
BRAM[3246]<= 32'hAAAAAAAA;
BRAM[3247]<= 32'hFFAAAAAA;
BRAM[3248]<= 32'hFFFFFFFF;
BRAM[3249]<= 32'hAAFEBFEA;
BRAM[3250]<= 32'hAAAAAAAA;
BRAM[3251]<= 32'hFAFFBFAA;
BRAM[3252]<= 32'hAAAAAAAA;
BRAM[3253]<= 32'hFAFFAFAA;
BRAM[3254]<= 32'hAAAAAAAA;
BRAM[3255]<= 32'hAAAAAAAA;
BRAM[3256]<= 32'hAAAAFFFF;
BRAM[3257]<= 32'hAAAAAAAA;
BRAM[3258]<= 32'hAAAAAAAA;
BRAM[3259]<= 32'hAAAAAAAA;
BRAM[3260]<= 32'hFFFFFFAF;
BRAM[3261]<= 32'hBFEAFFFF;
BRAM[3262]<= 32'hAAAAEAFF;
BRAM[3263]<= 32'hFFAAAAAA;
BRAM[3264]<= 32'hAAAAAAFF;
BRAM[3265]<= 32'hAAAAAAAA;
BRAM[3266]<= 32'hAAAAFFFF;
BRAM[3267]<= 32'hAAAAAAAA;
BRAM[3268]<= 32'hFEFFABAA;
BRAM[3269]<= 32'hAAAAAAAA;
BRAM[3270]<= 32'hAAAAAAAA;
BRAM[3271]<= 32'hAAAAAAAA;
BRAM[3272]<= 32'hFFFFAAAA;
BRAM[3273]<= 32'hFFFFFFFF;
BRAM[3274]<= 32'hFEFFBFEA;
BRAM[3275]<= 32'hAAAAAAAA;
BRAM[3276]<= 32'hAAFAFFAF;
BRAM[3277]<= 32'hAAAAAAAA;
BRAM[3278]<= 32'hFFAFAAAA;
BRAM[3279]<= 32'hAAAAAAFA;
BRAM[3280]<= 32'hBFAAAAAA;
BRAM[3281]<= 32'hAAAAEAFF;
BRAM[3282]<= 32'hAAAAAAAA;
BRAM[3283]<= 32'hAAAAAAAA;
BRAM[3284]<= 32'hAFAAAAAA;
BRAM[3285]<= 32'hFFFFFFFF;
BRAM[3286]<= 32'hBFEAFFFF;
BRAM[3287]<= 32'hAAEAFFFF;
BRAM[3288]<= 32'hFFFFAAAA;
BRAM[3289]<= 32'hAAAAAAAA;
BRAM[3290]<= 32'hAAAAAAAA;
BRAM[3291]<= 32'hAAFFFFAB;
BRAM[3292]<= 32'hAAAAAAAA;
BRAM[3293]<= 32'hAAFEFFAB;
BRAM[3294]<= 32'hAAAAAAAA;
BRAM[3295]<= 32'hAAAAAAAA;
BRAM[3296]<= 32'hAAAAAAAA;
BRAM[3297]<= 32'hFFFFFFAA;
BRAM[3298]<= 32'hFFFFFFFF;
BRAM[3299]<= 32'hFFFFBFEA;
BRAM[3300]<= 32'hAFAAAAFA;
BRAM[3301]<= 32'hAAAAFAFF;
BRAM[3302]<= 32'hAAAAAAAA;
BRAM[3303]<= 32'hBFAAAAAA;
BRAM[3304]<= 32'hAAAAEAFF;
BRAM[3305]<= 32'hFFBFAAAA;
BRAM[3306]<= 32'hAAAAAAEA;
BRAM[3307]<= 32'hAAAAAAAA;
BRAM[3308]<= 32'hAAAAAAAA;
BRAM[3309]<= 32'hFFABAAAA;
BRAM[3310]<= 32'hFFFFFFFF;
BRAM[3311]<= 32'hBFEAFFFF;
BRAM[3312]<= 32'hAAFFFFFF;
BRAM[3313]<= 32'hEAFFFFAA;
BRAM[3314]<= 32'hAAAAAAAA;
BRAM[3315]<= 32'hAAAAAAAA;
BRAM[3316]<= 32'hFEFFABAA;
BRAM[3317]<= 32'hABAAAAAA;
BRAM[3318]<= 32'hAAAAFEFF;
BRAM[3319]<= 32'hAAAAAAAA;
BRAM[3320]<= 32'hAAAAAAAA;
BRAM[3321]<= 32'hAAAAAAAA;
BRAM[3322]<= 32'hFFFFFFBF;
BRAM[3323]<= 32'hFFFFFFFF;
BRAM[3324]<= 32'hFFFFBFEA;
BRAM[3325]<= 32'hFFAFFAFF;
BRAM[3326]<= 32'hAAAAAAFE;
BRAM[3327]<= 32'hAAAAAAAA;
BRAM[3328]<= 32'hAAAAAAAA;
BRAM[3329]<= 32'hAAEAFFBF;
BRAM[3330]<= 32'hEAFFBFAA;
BRAM[3331]<= 32'hAAAAAAAA;
BRAM[3332]<= 32'hAAAAAAAA;
BRAM[3333]<= 32'hAAAAAAAA;
BRAM[3334]<= 32'hFFFFABAA;
BRAM[3335]<= 32'hFFFFFFFF;
BRAM[3336]<= 32'hBFEAFFFF;
BRAM[3337]<= 32'hFFFFFFFF;
BRAM[3338]<= 32'hAAEAFFBF;
BRAM[3339]<= 32'hAAAAAAAA;
BRAM[3340]<= 32'hAAAAAAAA;
BRAM[3341]<= 32'hFFABAAAA;
BRAM[3342]<= 32'hFFABAAFE;
BRAM[3343]<= 32'hAAAAAAFF;
BRAM[3344]<= 32'hAAAAAAAA;
BRAM[3345]<= 32'hAAAAAAAA;
BRAM[3346]<= 32'hBFAAAAAA;
BRAM[3347]<= 32'hFFFFFFFF;
BRAM[3348]<= 32'hFFFFFFFF;
BRAM[3349]<= 32'hFFFFBFEA;
BRAM[3350]<= 32'hFEFFFFFF;
BRAM[3351]<= 32'hAAAAAAAA;
BRAM[3352]<= 32'hAAAAAAAA;
BRAM[3353]<= 32'hAAAAAAAA;
BRAM[3354]<= 32'hAAFFFFAA;
BRAM[3355]<= 32'hAAFAFFAF;
BRAM[3356]<= 32'hAAAAAAAA;
BRAM[3357]<= 32'hAAAAAAAA;
BRAM[3358]<= 32'hAAAAAAAA;
BRAM[3359]<= 32'hFFFFFFAB;
BRAM[3360]<= 32'hFFFFFFFF;
BRAM[3361]<= 32'hBFEAFFFF;
BRAM[3362]<= 32'hFFFFFFFF;
BRAM[3363]<= 32'hAAAAEAFF;
BRAM[3364]<= 32'hAAAAAAAA;
BRAM[3365]<= 32'hAAAAAAAA;
BRAM[3366]<= 32'hAFAAAAAA;
BRAM[3367]<= 32'hFFFFFFFF;
BRAM[3368]<= 32'hAAAAAAAA;
BRAM[3369]<= 32'hAAAAAAAA;
BRAM[3370]<= 32'hAAAAAAAA;
BRAM[3371]<= 32'hFFBFAAAA;
BRAM[3372]<= 32'hFFFFFFFF;
BRAM[3373]<= 32'hFFFFFFFF;
BRAM[3374]<= 32'hFFFFBFEA;
BRAM[3375]<= 32'hEAFFFFFF;
BRAM[3376]<= 32'hAAAAAAAA;
BRAM[3377]<= 32'hAAAAAAAA;
BRAM[3378]<= 32'hAAAAAAAA;
BRAM[3379]<= 32'hFFFFAAAA;
BRAM[3380]<= 32'hAAAAFAFF;
BRAM[3381]<= 32'hAAAAAAAA;
BRAM[3382]<= 32'hAAAAAAAA;
BRAM[3383]<= 32'hABAAAAAA;
BRAM[3384]<= 32'hFFFFFFFF;
BRAM[3385]<= 32'hFFFFFFFF;
BRAM[3386]<= 32'hBFEAFFFF;
BRAM[3387]<= 32'hFFFFFFFF;
BRAM[3388]<= 32'hAAAAFEFF;
BRAM[3389]<= 32'hAAAAAAAA;
BRAM[3390]<= 32'hAAAAAAAA;
BRAM[3391]<= 32'hAAAAAAAA;
BRAM[3392]<= 32'hFAFFFFBF;
BRAM[3393]<= 32'hAAAAAAAA;
BRAM[3394]<= 32'hAAAAAAAA;
BRAM[3395]<= 32'hAAAAAAAA;
BRAM[3396]<= 32'hFFFFAFAA;
BRAM[3397]<= 32'hFFFFFFFF;
BRAM[3398]<= 32'hFFFFFFFF;
BRAM[3399]<= 32'hFFFFBFEA;
BRAM[3400]<= 32'hFFFFFFFF;
BRAM[3401]<= 32'hAAAAAAEA;
BRAM[3402]<= 32'hAAAAAAAA;
BRAM[3403]<= 32'hAAAAAAAA;
BRAM[3404]<= 32'hFFBFAAAA;
BRAM[3405]<= 32'hAAAAFAFF;
BRAM[3406]<= 32'hAAAAAAAA;
BRAM[3407]<= 32'hAAAAAAAA;
BRAM[3408]<= 32'hFFAAAAAA;
BRAM[3409]<= 32'hFFFFFFFF;
BRAM[3410]<= 32'hFFFFFFFF;
BRAM[3411]<= 32'hBFEAFFFF;
BRAM[3412]<= 32'hFFFFFFFF;
BRAM[3413]<= 32'hAAFAFFFF;
BRAM[3414]<= 32'hAAAAAAAA;
BRAM[3415]<= 32'hAAAAAAAA;
BRAM[3416]<= 32'hAAAAAAAA;
BRAM[3417]<= 32'hFAFFFFAF;
BRAM[3418]<= 32'hAAAAAAAA;
BRAM[3419]<= 32'hAAAAAAAA;
BRAM[3420]<= 32'hAAAAAAAA;
BRAM[3421]<= 32'hFFFFFFAF;
BRAM[3422]<= 32'hFFFFFFFF;
BRAM[3423]<= 32'hFFFFFFFF;
BRAM[3424]<= 32'hFFFFBFEA;
BRAM[3425]<= 32'hFFFFFFFF;
BRAM[3426]<= 32'hAAAAAAFF;
BRAM[3427]<= 32'hAAAAAAAA;
BRAM[3428]<= 32'hAAAAAAAA;
BRAM[3429]<= 32'hFFABAAAA;
BRAM[3430]<= 32'hAAAAFEFF;
BRAM[3431]<= 32'hAAAAAAAA;
BRAM[3432]<= 32'hAAAAAAAA;
BRAM[3433]<= 32'hFFFFAAAA;
BRAM[3434]<= 32'hFFFFFFFF;
BRAM[3435]<= 32'hFFFFFFFF;
BRAM[3436]<= 32'hBFEAFFFF;
BRAM[3437]<= 32'hFFFFFFFF;
BRAM[3438]<= 32'hFAFFFFFF;
BRAM[3439]<= 32'hAAAAAAAA;
BRAM[3440]<= 32'hAAAAAAAA;
BRAM[3441]<= 32'hAAAAAAAA;
BRAM[3442]<= 32'hFFFFBFAA;
BRAM[3443]<= 32'hAAAAAAEA;
BRAM[3444]<= 32'hAAAAAAAA;
BRAM[3445]<= 32'hAFAAAAAA;
BRAM[3446]<= 32'hFFFFFFFF;
BRAM[3447]<= 32'hFFFFFFFF;
BRAM[3448]<= 32'hFFFFFFFF;
BRAM[3449]<= 32'hFFFFBFEA;
BRAM[3450]<= 32'hFFFFFFFF;
BRAM[3451]<= 32'hAAAAFFFF;
BRAM[3452]<= 32'hAAAAAAAA;
BRAM[3453]<= 32'hAAAAAAAA;
BRAM[3454]<= 32'hAAAAAAAA;
BRAM[3455]<= 32'hAAFEFFAB;
BRAM[3456]<= 32'hAAAAAAAA;
BRAM[3457]<= 32'hAAAAAAAA;
BRAM[3458]<= 32'hFFFFFFAA;
BRAM[3459]<= 32'hFFFFFFFF;
BRAM[3460]<= 32'hFFFFFFFF;
BRAM[3461]<= 32'hBFEAFFFF;
BRAM[3462]<= 32'hFFFFFFFF;
BRAM[3463]<= 32'hFFFFFFFF;
BRAM[3464]<= 32'hAAAAAAEA;
BRAM[3465]<= 32'hAAAAAAAA;
BRAM[3466]<= 32'hAAAAAAAA;
BRAM[3467]<= 32'hFFAAAAAA;
BRAM[3468]<= 32'hAAAAAAFF;
BRAM[3469]<= 32'hAAAAAAAA;
BRAM[3470]<= 32'hFFAFAAAA;
BRAM[3471]<= 32'hFFFFFFFF;
BRAM[3472]<= 32'hFFFFFFFF;
BRAM[3473]<= 32'hFFFFFFFF;
BRAM[3474]<= 32'hFFFFBFEA;
BRAM[3475]<= 32'hFFFFFFFF;
BRAM[3476]<= 32'hAAFEFFFF;
BRAM[3477]<= 32'hAAAAAAAA;
BRAM[3478]<= 32'hAAAAAAAA;
BRAM[3479]<= 32'hAAAAAAAA;
BRAM[3480]<= 32'hFAFFAFAA;
BRAM[3481]<= 32'hAAAAAAAA;
BRAM[3482]<= 32'hAAAAAAAA;
BRAM[3483]<= 32'hFFFFFFBF;
BRAM[3484]<= 32'hFFFFFFF6;
BRAM[3485]<= 32'hFFFFFFFF;
BRAM[3486]<= 32'hBFEAFFFF;
BRAM[3487]<= 32'hFFFFFFFF;
BRAM[3488]<= 32'hFFFFFFFF;
BRAM[3489]<= 32'hAAAAEAFF;
BRAM[3490]<= 32'hAAAAAAAA;
BRAM[3491]<= 32'hAAAAAAAA;
BRAM[3492]<= 32'hAAAAAAAA;
BRAM[3493]<= 32'hAAAAFFFF;
BRAM[3494]<= 32'hAAAAAAAA;
BRAM[3495]<= 32'hFFFFABAA;
BRAM[3496]<= 32'hFF81FFFF;
BRAM[3497]<= 32'hFFFFFFFF;
BRAM[3498]<= 32'hFFFFFFFF;
BRAM[3499]<= 32'hFFFFBFEA;
BRAM[3500]<= 32'hBFFFFFFF;
BRAM[3501]<= 32'hFEFFFFFF;
BRAM[3502]<= 32'hAAAAAAAA;
BRAM[3503]<= 32'hAAAAAAAA;
BRAM[3504]<= 32'hAAAAAAAA;
BRAM[3505]<= 32'hFFAFAAAA;
BRAM[3506]<= 32'hAAAAAAFA;
BRAM[3507]<= 32'hBFAAAAAA;
BRAM[3508]<= 32'hF8FFFFFF;
BRAM[3509]<= 32'hFFFFFF00;
BRAM[3510]<= 32'hFFFFFFFF;
BRAM[3511]<= 32'hBFEAFFFF;
BRAM[3512]<= 32'hFFFFFFFF;
BRAM[3513]<= 32'hFFFF07FF;
BRAM[3514]<= 32'hAAEAFFFF;
BRAM[3515]<= 32'hAAAAAAAA;
BRAM[3516]<= 32'hAAAAAAAA;
BRAM[3517]<= 32'hAAAAAAAA;
BRAM[3518]<= 32'hAAFFFFAB;
BRAM[3519]<= 32'hAAAAAAAA;
BRAM[3520]<= 32'hFFFFFFAB;
BRAM[3521]<= 32'hBF00D0FF;
BRAM[3522]<= 32'hFFFFFFFF;
BRAM[3523]<= 32'hFFFFFFFF;
BRAM[3524]<= 32'hFFFFBFEA;
BRAM[3525]<= 32'h00FEFFFF;
BRAM[3526]<= 32'hFFFFFFBF;
BRAM[3527]<= 32'hAAAAAAFA;
BRAM[3528]<= 32'hAAAAAAAA;
BRAM[3529]<= 32'hAAAAAAAA;
BRAM[3530]<= 32'hBFAAAAAA;
BRAM[3531]<= 32'hAAAAEAFF;
BRAM[3532]<= 32'hFFBFAAAA;
BRAM[3533]<= 32'h00FDFFFF;
BRAM[3534]<= 32'hFFFF7F00;
BRAM[3535]<= 32'hFFFFFFFF;
BRAM[3536]<= 32'hBFEAFFFF;
BRAM[3537]<= 32'hFFFFFFFF;
BRAM[3538]<= 32'hFF0B00FD;
BRAM[3539]<= 32'hAAFFFFFF;
BRAM[3540]<= 32'hAAAAAAAA;
BRAM[3541]<= 32'hAAAAAAAA;
BRAM[3542]<= 32'hAAAAAAAA;
BRAM[3543]<= 32'hFEFFABAA;
BRAM[3544]<= 32'hABAAAAAA;
BRAM[3545]<= 32'hFFFFFFFF;
BRAM[3546]<= 32'h3F0000E0;
BRAM[3547]<= 32'hFFFFFFFF;
BRAM[3548]<= 32'hFFFFFFFF;
BRAM[3549]<= 32'hFFFFBFEA;
BRAM[3550]<= 32'h00FCFFFF;
BRAM[3551]<= 32'hFFFFBF01;
BRAM[3552]<= 32'hAAAAFAFF;
BRAM[3553]<= 32'hAAAAAAAA;
BRAM[3554]<= 32'hAAAAAAAA;
BRAM[3555]<= 32'hAAAAAAAA;
BRAM[3556]<= 32'hAAEAFFBF;
BRAM[3557]<= 32'hFFFFBFAA;
BRAM[3558]<= 32'h0000FEFF;
BRAM[3559]<= 32'hFFFF3F00;
BRAM[3560]<= 32'hFFFFFFFF;
BRAM[3561]<= 32'hBFEAFFFF;
BRAM[3562]<= 32'hFFFFFFFF;
BRAM[3563]<= 32'h1F0000FC;
BRAM[3564]<= 32'hFFFFFFFF;
BRAM[3565]<= 32'hAAAAAAAA;
BRAM[3566]<= 32'hAAAAAAAA;
BRAM[3567]<= 32'hAAAAAAAA;
BRAM[3568]<= 32'hFFABAAAA;
BRAM[3569]<= 32'hFFAAAAFE;
BRAM[3570]<= 32'hE4FFFFFF;
BRAM[3571]<= 32'h2F000000;
BRAM[3572]<= 32'hFFFFFFFF;
BRAM[3573]<= 32'hFEFFFFFF;
BRAM[3574]<= 32'hFFFFABAA;
BRAM[3575]<= 32'h00F8FFFF;
BRAM[3576]<= 32'hFFFF0100;
BRAM[3577]<= 32'hAAFAFFFF;
BRAM[3578]<= 32'hAAAAAAAA;
BRAM[3579]<= 32'hAAAAAAAA;
BRAM[3580]<= 32'hAAAAAAAA;
BRAM[3581]<= 32'hAAFFFFAA;
BRAM[3582]<= 32'hFFFFFFAF;
BRAM[3583]<= 32'h000040FF;
BRAM[3584]<= 32'hFFFF1F00;
BRAM[3585]<= 32'hFFFFFFFF;
BRAM[3586]<= 32'hAAAAFAFF;
BRAM[3587]<= 32'hFFFFFFFF;
BRAM[3588]<= 32'h000000F4;
BRAM[3589]<= 32'hFFFFFF2F;
BRAM[3590]<= 32'hAAAAAAFE;
BRAM[3591]<= 32'hAAAAAAAA;
BRAM[3592]<= 32'hAAAAAAAA;
BRAM[3593]<= 32'hAFAAAAAA;
BRAM[3594]<= 32'hFFFFFAFF;
BRAM[3595]<= 32'h00F4FFFF;
BRAM[3596]<= 32'h0F000000;
BRAM[3597]<= 32'hFFFFFFFF;
BRAM[3598]<= 32'hFAFFFFFF;
BRAM[3599]<= 32'hFFFFAAAA;
BRAM[3600]<= 32'h00F0FFFF;
BRAM[3601]<= 32'hFF020000;
BRAM[3602]<= 32'hEAFFFFFF;
BRAM[3603]<= 32'hAAAAAAAA;
BRAM[3604]<= 32'hAAAAAAAA;
BRAM[3605]<= 32'hAAAAAAAA;
BRAM[3606]<= 32'hFFFFAAAA;
BRAM[3607]<= 32'hFFFFFFFF;
BRAM[3608]<= 32'h00000080;
BRAM[3609]<= 32'hFFFF0F00;
BRAM[3610]<= 32'hFFFFFFFF;
BRAM[3611]<= 32'hAAAAEAFF;
BRAM[3612]<= 32'hFFFFFFBF;
BRAM[3613]<= 32'h000000F0;
BRAM[3614]<= 32'hFFFF7F00;
BRAM[3615]<= 32'hAAAAFEFF;
BRAM[3616]<= 32'hAAAAAAAA;
BRAM[3617]<= 32'hAAAAAAAA;
BRAM[3618]<= 32'hAAAAAAAA;
BRAM[3619]<= 32'hFFFFFFAF;
BRAM[3620]<= 32'h0000F8FF;
BRAM[3621]<= 32'h0B000000;
BRAM[3622]<= 32'hFFFFFFFF;
BRAM[3623]<= 32'hEAFFFFFF;
BRAM[3624]<= 32'hFFBFAAAA;
BRAM[3625]<= 32'h00E0FFFF;
BRAM[3626]<= 32'h07000000;
BRAM[3627]<= 32'hFFFFFFFF;
BRAM[3628]<= 32'hAAAAAAEA;
BRAM[3629]<= 32'hAAAAAAAA;
BRAM[3630]<= 32'hAAAAAAAA;
BRAM[3631]<= 32'hFFAFAAAA;
BRAM[3632]<= 32'h90FFFFFF;
BRAM[3633]<= 32'h00000000;
BRAM[3634]<= 32'hFFFF0B00;
BRAM[3635]<= 32'hFFFFFFFF;
BRAM[3636]<= 32'hAAAAEAFF;
BRAM[3637]<= 32'hFFFFFFBF;
BRAM[3638]<= 32'h000000D0;
BRAM[3639]<= 32'hFFBF0000;
BRAM[3640]<= 32'hAAFAFFFF;
BRAM[3641]<= 32'hAAAAAAAA;
BRAM[3642]<= 32'hAAAAAAAA;
BRAM[3643]<= 32'hAAAAAAAA;
BRAM[3644]<= 32'hFFFFFFFF;
BRAM[3645]<= 32'h000000FD;
BRAM[3646]<= 32'h07000000;
BRAM[3647]<= 32'hFFFFFFFF;
BRAM[3648]<= 32'hEAFFFFFF;
BRAM[3649]<= 32'hFFBFAAAA;
BRAM[3650]<= 32'h00D0FFFF;
BRAM[3651]<= 32'h00000000;
BRAM[3652]<= 32'hFFFFFF0B;
BRAM[3653]<= 32'hAAAAAAFF;
BRAM[3654]<= 32'hAAAAAAAA;
BRAM[3655]<= 32'hAAAAAAAA;
BRAM[3656]<= 32'hFFFFABAA;
BRAM[3657]<= 32'h00D0FFFF;
BRAM[3658]<= 32'h00000000;
BRAM[3659]<= 32'hFFFF0300;
BRAM[3660]<= 32'hFFFFFFFF;
BRAM[3661]<= 32'hAAAAEAFF;
BRAM[3662]<= 32'hFFFFFFBF;
BRAM[3663]<= 32'h000000C0;
BRAM[3664]<= 32'hBF010000;
BRAM[3665]<= 32'hFAFFFFFF;
BRAM[3666]<= 32'hAAAAAAAA;
BRAM[3667]<= 32'hAAAAAAAA;
BRAM[3668]<= 32'hBFAAAAAA;
BRAM[3669]<= 32'hFEFFFFFF;
BRAM[3670]<= 32'h00000000;
BRAM[3671]<= 32'h03000000;
BRAM[3672]<= 32'hFFFFFFFF;
BRAM[3673]<= 32'hEAFFFFFF;
BRAM[3674]<= 32'hFFBFAAAA;
BRAM[3675]<= 32'h00C0FFFF;
BRAM[3676]<= 32'h00000000;
BRAM[3677]<= 32'hFFFF1F00;
BRAM[3678]<= 32'hAAAAFFFF;
BRAM[3679]<= 32'hAAAAAAAA;
BRAM[3680]<= 32'hAAAAAAAA;
BRAM[3681]<= 32'hFFFFFFAB;
BRAM[3682]<= 32'h0000E0FF;
BRAM[3683]<= 32'h00000000;
BRAM[3684]<= 32'hFFFF0200;
BRAM[3685]<= 32'hFFFFFFFF;
BRAM[3686]<= 32'hAAAAEAFF;
BRAM[3687]<= 32'hFFFFFFBF;
BRAM[3688]<= 32'h00000080;
BRAM[3689]<= 32'h01000000;
BRAM[3690]<= 32'hFFFFFFFF;
BRAM[3691]<= 32'hAAAAAAFA;
BRAM[3692]<= 32'hAAAAAAAA;
BRAM[3693]<= 32'hFFBFAAAA;
BRAM[3694]<= 32'h40FEFFFF;
BRAM[3695]<= 32'h00000000;
BRAM[3696]<= 32'h01000000;
BRAM[3697]<= 32'hFFFFFFFF;
BRAM[3698]<= 32'hEAFFFFFF;
BRAM[3699]<= 32'hFFBFAAAA;
BRAM[3700]<= 32'h0040FFFF;
BRAM[3701]<= 32'h00000000;
BRAM[3702]<= 32'hFF2F0000;
BRAM[3703]<= 32'hAAFEFFFF;
BRAM[3704]<= 32'hAAAAAAAA;
BRAM[3705]<= 32'hABAAAAAA;
BRAM[3706]<= 32'hFFFFFFFF;
BRAM[3707]<= 32'h000000F4;
BRAM[3708]<= 32'h00000000;
BRAM[3709]<= 32'hFFFF0100;
BRAM[3710]<= 32'hFFFFFFFF;
BRAM[3711]<= 32'hAAAAEAFF;
BRAM[3712]<= 32'hFFFFFFBF;
BRAM[3713]<= 32'h00000040;
BRAM[3714]<= 32'h00000000;
BRAM[3715]<= 32'hFFFFFF02;
BRAM[3716]<= 32'hAAAAEAFF;
BRAM[3717]<= 32'hAAAAAAAA;
BRAM[3718]<= 32'hFFFFBFAA;
BRAM[3719]<= 32'h0040FFFF;
BRAM[3720]<= 32'h00000000;
BRAM[3721]<= 32'h00000000;
BRAM[3722]<= 32'hFFFFFFFF;
BRAM[3723]<= 32'hEAFFFFFF;
BRAM[3724]<= 32'hFFBFAAAA;
BRAM[3725]<= 32'h0000FFFF;
BRAM[3726]<= 32'h00000000;
BRAM[3727]<= 32'h7F000000;
BRAM[3728]<= 32'hFEFFFFFF;
BRAM[3729]<= 32'hAAAAAAAA;
BRAM[3730]<= 32'hFFABAAAA;
BRAM[3731]<= 32'hF4FFFFFF;
BRAM[3732]<= 32'h00000000;
BRAM[3733]<= 32'h00000000;
BRAM[3734]<= 32'hFFFF0000;
BRAM[3735]<= 32'hFFFFFFFF;
BRAM[3736]<= 32'hAAAAEAFF;
BRAM[3737]<= 32'hFFFFFFBF;
BRAM[3738]<= 32'h00000000;
BRAM[3739]<= 32'h00000000;
BRAM[3740]<= 32'hFFFF0700;
BRAM[3741]<= 32'hAAEAFFFF;
BRAM[3742]<= 32'hAAAAAAAA;
BRAM[3743]<= 32'hFFFFFFAF;
BRAM[3744]<= 32'h000080FF;
BRAM[3745]<= 32'h00000000;
BRAM[3746]<= 32'h00000000;
BRAM[3747]<= 32'hFFFFFFBF;
BRAM[3748]<= 32'hEAFFFFFF;
BRAM[3749]<= 32'hFFBFAAAA;
BRAM[3750]<= 32'h0000FEFF;
BRAM[3751]<= 32'h00000000;
BRAM[3752]<= 32'h00000000;
BRAM[3753]<= 32'hFFFFFFBF;
BRAM[3754]<= 32'hAAAAAAFA;
BRAM[3755]<= 32'hFFFFAAAA;
BRAM[3756]<= 32'h00F8FFFF;
BRAM[3757]<= 32'h00000000;
BRAM[3758]<= 32'h00000000;
BRAM[3759]<= 32'hFF7F0000;
BRAM[3760]<= 32'hFFFFFFFF;
BRAM[3761]<= 32'hAAAAEAFF;
BRAM[3762]<= 32'hFDFFFFBF;
BRAM[3763]<= 32'h00000000;
BRAM[3764]<= 32'h00000000;
BRAM[3765]<= 32'hFF0B0000;
BRAM[3766]<= 32'hAAFFFFFF;
BRAM[3767]<= 32'hAFAAAAAA;
BRAM[3768]<= 32'hFFFFFFFF;
BRAM[3769]<= 32'h00000090;
BRAM[3770]<= 32'h00000000;
BRAM[3771]<= 32'h00000000;
BRAM[3772]<= 32'hFFFFFF7F;
BRAM[3773]<= 32'hEAFFFFFF;
BRAM[3774]<= 32'hFFBFAAAA;
BRAM[3775]<= 32'h0000FDFF;
BRAM[3776]<= 32'h00000000;
BRAM[3777]<= 32'h00000000;
BRAM[3778]<= 32'hFFFFBF00;
BRAM[3779]<= 32'hAAAAFAFF;
BRAM[3780]<= 32'hFFFFFFAA;
BRAM[3781]<= 32'h0000FDFF;
BRAM[3782]<= 32'h00000000;
BRAM[3783]<= 32'h00000000;
BRAM[3784]<= 32'hFF3F0000;
BRAM[3785]<= 32'hFFFFFFFF;
BRAM[3786]<= 32'hAAAAEAFF;
BRAM[3787]<= 32'hFCFFFFBF;
BRAM[3788]<= 32'h00000000;
BRAM[3789]<= 32'h00000000;
BRAM[3790]<= 32'h1F000000;
BRAM[3791]<= 32'hFFFFFFFF;
BRAM[3792]<= 32'hFFAFAAAA;
BRAM[3793]<= 32'hD0FFFFFF;
BRAM[3794]<= 32'h00000000;
BRAM[3795]<= 32'h00000000;
BRAM[3796]<= 32'h00000000;
BRAM[3797]<= 32'hFFFFFF3F;
BRAM[3798]<= 32'hEAFFFFFF;
BRAM[3799]<= 32'hFFBFAAAA;
BRAM[3800]<= 32'h0000FCFF;
BRAM[3801]<= 32'h00000000;
BRAM[3802]<= 32'h00000000;
BRAM[3803]<= 32'hFFFF0100;
BRAM[3804]<= 32'hFFFFFFFF;
BRAM[3805]<= 32'hFFFFFFFF;
BRAM[3806]<= 32'h000000FD;
BRAM[3807]<= 32'h00000000;
BRAM[3808]<= 32'h00000000;
BRAM[3809]<= 32'hFF3F0000;
BRAM[3810]<= 32'hFFFFFFFF;
BRAM[3811]<= 32'hAAAAEAFF;
BRAM[3812]<= 32'hFCFFFFBF;
BRAM[3813]<= 32'h00000000;
BRAM[3814]<= 32'h00000000;
BRAM[3815]<= 32'h00000000;
BRAM[3816]<= 32'hFFFFFF2F;
BRAM[3817]<= 32'hFFFFFFFF;
BRAM[3818]<= 32'h00E0FFFF;
BRAM[3819]<= 32'h00000000;
BRAM[3820]<= 32'h00000000;
BRAM[3821]<= 32'h00000000;
BRAM[3822]<= 32'hFFFFFF2F;
BRAM[3823]<= 32'hEAFFFFFF;
BRAM[3824]<= 32'hFFBFAAAA;
BRAM[3825]<= 32'h0000F8FF;
BRAM[3826]<= 32'h00000000;
BRAM[3827]<= 32'h00000000;
BRAM[3828]<= 32'hFF020000;
BRAM[3829]<= 32'hFFFFFFFF;
BRAM[3830]<= 32'hFEFFFFFF;
BRAM[3831]<= 32'h00000000;
BRAM[3832]<= 32'h00000000;
BRAM[3833]<= 32'h00000000;
BRAM[3834]<= 32'hFF2F0000;
BRAM[3835]<= 32'hFFFFFFFF;
BRAM[3836]<= 32'hAAAAEAFF;
BRAM[3837]<= 32'hF8FFFFBF;
BRAM[3838]<= 32'h00000000;
BRAM[3839]<= 32'h00000000;
BRAM[3840]<= 32'h00000000;
BRAM[3841]<= 32'hFFFF6F00;
BRAM[3842]<= 32'hFFFFFFFF;
BRAM[3843]<= 32'h0000E4FF;
BRAM[3844]<= 32'h00000000;
BRAM[3845]<= 32'h00000000;
BRAM[3846]<= 32'h00000000;
BRAM[3847]<= 32'hFFFFFF1F;
BRAM[3848]<= 32'hEAFFFFFF;
BRAM[3849]<= 32'hFFBFAAAA;
BRAM[3850]<= 32'h0000F8FF;
BRAM[3851]<= 32'h00000000;
BRAM[3852]<= 32'h00000000;
BRAM[3853]<= 32'h07000000;
BRAM[3854]<= 32'hFFFFFFFF;
BRAM[3855]<= 32'h40FFFFFF;
BRAM[3856]<= 32'h00000000;
BRAM[3857]<= 32'h00000000;
BRAM[3858]<= 32'h00000000;
BRAM[3859]<= 32'hFF1F0000;
BRAM[3860]<= 32'hFFFFFFFF;
BRAM[3861]<= 32'hAAAAEAFF;
BRAM[3862]<= 32'hF4FFFFBF;
BRAM[3863]<= 32'h00000000;
BRAM[3864]<= 32'h00000000;
BRAM[3865]<= 32'h00000000;
BRAM[3866]<= 32'hFF7F0000;
BRAM[3867]<= 32'hFFFFFFFF;
BRAM[3868]<= 32'h000000F4;
BRAM[3869]<= 32'h00000000;
BRAM[3870]<= 32'h00000000;
BRAM[3871]<= 32'h00000000;
BRAM[3872]<= 32'hFFFFFF1F;
BRAM[3873]<= 32'hEAFFFFFF;
BRAM[3874]<= 32'hFFBFAAAA;
BRAM[3875]<= 32'h0000F4FF;
BRAM[3876]<= 32'h00000000;
BRAM[3877]<= 32'h00000000;
BRAM[3878]<= 32'h00000000;
BRAM[3879]<= 32'hFFFFFF0B;
BRAM[3880]<= 32'h0080FFFF;
BRAM[3881]<= 32'h00000000;
BRAM[3882]<= 32'h00000000;
BRAM[3883]<= 32'h00000000;
BRAM[3884]<= 32'hFF1F0000;
BRAM[3885]<= 32'hFFFFFFFF;
BRAM[3886]<= 32'hAAAAEAFF;
BRAM[3887]<= 32'hF4FFFFBF;
BRAM[3888]<= 32'h00000000;
BRAM[3889]<= 32'h00000000;
BRAM[3890]<= 32'h00000000;
BRAM[3891]<= 32'hBF000000;
BRAM[3892]<= 32'hF8FFFFFF;
BRAM[3893]<= 32'h00000000;
BRAM[3894]<= 32'h00000000;
BRAM[3895]<= 32'h00000000;
BRAM[3896]<= 32'h00000000;
BRAM[3897]<= 32'hFFFFFF0F;
BRAM[3898]<= 32'hEAFFFFFF;
BRAM[3899]<= 32'hFFBFAAAA;
BRAM[3900]<= 32'h0000F8FF;
BRAM[3901]<= 32'h00000000;
BRAM[3902]<= 32'h00000000;
BRAM[3903]<= 32'h00000000;
BRAM[3904]<= 32'hFFFF1F00;
BRAM[3905]<= 32'h0000D0FF;
BRAM[3906]<= 32'h00000000;
BRAM[3907]<= 32'h00000000;
BRAM[3908]<= 32'h00000000;
BRAM[3909]<= 32'hFF2F0000;
BRAM[3910]<= 32'hFFFFFFFF;
BRAM[3911]<= 32'hAAAAEAFF;
BRAM[3912]<= 32'hFFFFFFBF;
BRAM[3913]<= 32'h000000F9;
BRAM[3914]<= 32'h00000000;
BRAM[3915]<= 32'h00000000;
BRAM[3916]<= 32'h01000000;
BRAM[3917]<= 32'h00FEFFFF;
BRAM[3918]<= 32'h00000000;
BRAM[3919]<= 32'h00000000;
BRAM[3920]<= 32'h00000000;
BRAM[3921]<= 32'h6F000000;
BRAM[3922]<= 32'hFFFFFFFF;
BRAM[3923]<= 32'hEAFFFFFF;
BRAM[3924]<= 32'hFFBFAAAA;
BRAM[3925]<= 32'hF9FFFFFF;
BRAM[3926]<= 32'h00000000;
BRAM[3927]<= 32'h00000000;
BRAM[3928]<= 32'h00000000;
BRAM[3929]<= 32'hFF0A0000;
BRAM[3930]<= 32'h000000E0;
BRAM[3931]<= 32'h00000000;
BRAM[3932]<= 32'h00000000;
BRAM[3933]<= 32'h00000000;
BRAM[3934]<= 32'hFFFFFF6F;
BRAM[3935]<= 32'hFFFFFFFF;
BRAM[3936]<= 32'hAAAAEAFF;
BRAM[3937]<= 32'hFFFFFFBF;
BRAM[3938]<= 32'h00E4FFFF;
BRAM[3939]<= 32'h00000000;
BRAM[3940]<= 32'h00000000;
BRAM[3941]<= 32'h00000000;
BRAM[3942]<= 32'h00000000;
BRAM[3943]<= 32'h00000000;
BRAM[3944]<= 32'h00000000;
BRAM[3945]<= 32'h00000000;
BRAM[3946]<= 32'hFFFF1B00;
BRAM[3947]<= 32'hFFFFFFFF;
BRAM[3948]<= 32'hEAFFFFFF;
BRAM[3949]<= 32'hFFBFAAAA;
BRAM[3950]<= 32'hFFFFFFFF;
BRAM[3951]<= 32'h0000D0FF;
BRAM[3952]<= 32'h00000000;
BRAM[3953]<= 32'h00000000;
BRAM[3954]<= 32'h00000000;
BRAM[3955]<= 32'h00000000;
BRAM[3956]<= 32'h00000000;
BRAM[3957]<= 32'h00000000;
BRAM[3958]<= 32'hFF060000;
BRAM[3959]<= 32'hFFFFFFFF;
BRAM[3960]<= 32'hFFFFFFFF;
BRAM[3961]<= 32'hAAAAAAFF;
BRAM[3962]<= 32'hFFFFFFBF;
BRAM[3963]<= 32'hFFFFFFFF;
BRAM[3964]<= 32'h00000080;
BRAM[3965]<= 32'h00000000;
BRAM[3966]<= 32'h00000000;
BRAM[3967]<= 32'h00000000;
BRAM[3968]<= 32'h00000000;
BRAM[3969]<= 32'h00000000;
BRAM[3970]<= 32'h01000000;
BRAM[3971]<= 32'hFFFFFFBF;
BRAM[3972]<= 32'hFFFFFFFF;
BRAM[3973]<= 32'hAAFFFFFF;
BRAM[3974]<= 32'hFFBFAEAA;
BRAM[3975]<= 32'hFFFFFFFF;
BRAM[3976]<= 32'h00FDFFFF;
BRAM[3977]<= 32'h00000000;
BRAM[3978]<= 32'h00000000;
BRAM[3979]<= 32'h00000000;
BRAM[3980]<= 32'h00000000;
BRAM[3981]<= 32'h00000000;
BRAM[3982]<= 32'h00000000;
BRAM[3983]<= 32'hFFFF6F00;
BRAM[3984]<= 32'hFFFFFFFF;
BRAM[3985]<= 32'hFFFFFFFF;
BRAM[3986]<= 32'hFFBAABFF;
BRAM[3987]<= 32'hFFFFFFBF;
BRAM[3988]<= 32'hFFFFFFFF;
BRAM[3989]<= 32'h0000E4FF;
BRAM[3990]<= 32'h00000000;
BRAM[3991]<= 32'h00000000;
BRAM[3992]<= 32'h00000000;
BRAM[3993]<= 32'h00000000;
BRAM[3994]<= 32'h00000000;
BRAM[3995]<= 32'hFF1B0000;
BRAM[3996]<= 32'hFFFFFFFF;
BRAM[3997]<= 32'hFFFFFFFF;
BRAM[3998]<= 32'hABFFFFFF;
BRAM[3999]<= 32'hFFBFFFBA;
BRAM[4000]<= 32'hFFFFFFFF;
BRAM[4001]<= 32'hFFFFFFFF;
BRAM[4002]<= 32'h00000090;
BRAM[4003]<= 32'h00000000;
BRAM[4004]<= 32'h00000000;
BRAM[4005]<= 32'h00000000;
BRAM[4006]<= 32'h00000000;
BRAM[4007]<= 32'h06000000;
BRAM[4008]<= 32'hFFFFFFFF;
BRAM[4009]<= 32'hFFFFFFFF;
BRAM[4010]<= 32'hFFFFFFFF;
BRAM[4011]<= 32'hFFBAABFF;
BRAM[4012]<= 32'hFFFFFFBF;
BRAM[4013]<= 32'hFFFFFFFF;
BRAM[4014]<= 32'h00FEFFFF;
BRAM[4015]<= 32'h00000000;
BRAM[4016]<= 32'h00000000;
BRAM[4017]<= 32'h00000000;
BRAM[4018]<= 32'h00000000;
BRAM[4019]<= 32'h00000000;
BRAM[4020]<= 32'hFFFF7F00;
BRAM[4021]<= 32'hFFFFFFFF;
BRAM[4022]<= 32'hFFFFFFFF;
BRAM[4023]<= 32'hABFFFFFF;
BRAM[4024]<= 32'hFFBFFFBA;
BRAM[4025]<= 32'hFFFFFFFF;
BRAM[4026]<= 32'hFFFFFFFF;
BRAM[4027]<= 32'h0000F4FF;
BRAM[4028]<= 32'h00000000;
BRAM[4029]<= 32'h00000000;
BRAM[4030]<= 32'h00000000;
BRAM[4031]<= 32'h00000000;
BRAM[4032]<= 32'hFF1B0000;
BRAM[4033]<= 32'hFFFFFFFF;
BRAM[4034]<= 32'hFFFFFFFF;
BRAM[4035]<= 32'hFFFFFFFF;
BRAM[4036]<= 32'hFFBAABFF;
BRAM[4037]<= 32'hFFFFFFBF;
BRAM[4038]<= 32'hFFFFFFFF;
BRAM[4039]<= 32'hFFFFFFFF;
BRAM[4040]<= 32'h00000080;
BRAM[4041]<= 32'h00000000;
BRAM[4042]<= 32'h00000000;
BRAM[4043]<= 32'h00000000;
BRAM[4044]<= 32'h02000000;
BRAM[4045]<= 32'hFFFFFFFF;
BRAM[4046]<= 32'hFFFFFFFF;
BRAM[4047]<= 32'hFFFFFFFF;
BRAM[4048]<= 32'hABFFFFFF;
BRAM[4049]<= 32'hFFBFFFBA;
BRAM[4050]<= 32'hFFFFFFFF;
BRAM[4051]<= 32'hFFFFFFFF;
BRAM[4052]<= 32'h00F9FFFF;
BRAM[4053]<= 32'h00000000;
BRAM[4054]<= 32'h00000000;
BRAM[4055]<= 32'h00000000;
BRAM[4056]<= 32'h00000000;
BRAM[4057]<= 32'hFFFF6F00;
BRAM[4058]<= 32'hFFFFFFFF;
BRAM[4059]<= 32'hFFFFFFFF;
BRAM[4060]<= 32'hFFFFFFFF;
BRAM[4061]<= 32'hFFBAABFF;
BRAM[4062]<= 32'hFFFFFFBF;
BRAM[4063]<= 32'hFFFFFFFF;
BRAM[4064]<= 32'hFFFFFFFF;
BRAM[4065]<= 32'h0000D0FF;
BRAM[4066]<= 32'h00000000;
BRAM[4067]<= 32'h00000000;
BRAM[4068]<= 32'h00000000;
BRAM[4069]<= 32'hFF070000;
BRAM[4070]<= 32'hFFFFFFFF;
BRAM[4071]<= 32'hFFFFFFFF;
BRAM[4072]<= 32'hFFFFFFFF;
BRAM[4073]<= 32'hABFFFFFF;
BRAM[4074]<= 32'hFFBFFFBA;
BRAM[4075]<= 32'hFFFFFFFF;
BRAM[4076]<= 32'hFFFFFFFF;
BRAM[4077]<= 32'hFEFFFFFF;
BRAM[4078]<= 32'h00000000;
BRAM[4079]<= 32'h00000000;
BRAM[4080]<= 32'h00000000;
BRAM[4081]<= 32'h00000000;
BRAM[4082]<= 32'hFFFFFFBF;
BRAM[4083]<= 32'hFFFFFFFF;
BRAM[4084]<= 32'hFFFFFFFF;
BRAM[4085]<= 32'hFFFFFFFF;
BRAM[4086]<= 32'hFFBAABFF;
BRAM[4087]<= 32'hFFFFFFBF;
BRAM[4088]<= 32'hFFFFFFFF;
BRAM[4089]<= 32'hFFFFFFFF;
BRAM[4090]<= 32'h00E4FFFF;
BRAM[4091]<= 32'h00000000;
BRAM[4092]<= 32'h00000000;
BRAM[4093]<= 32'h00000000;
BRAM[4094]<= 32'hFFFF0B00;
BRAM[4095]<= 32'hFFFFFFFF;
BRAM[4096]<= 32'hFFFFFFFF;
BRAM[4097]<= 32'hFFFFFFFF;
BRAM[4098]<= 32'hABFFFFFF;
BRAM[4099]<= 32'hFFBFFFBA;
BRAM[4100]<= 32'hFFFFFFFF;
BRAM[4101]<= 32'hFFFFFFFF;
BRAM[4102]<= 32'hFFFFFFFF;
BRAM[4103]<= 32'h000040FF;
BRAM[4104]<= 32'h00000000;
BRAM[4105]<= 32'h00000000;
BRAM[4106]<= 32'hBF010000;
BRAM[4107]<= 32'hFFFFFFFF;
BRAM[4108]<= 32'hFFFFFFFF;
BRAM[4109]<= 32'hFFFFFFFF;
BRAM[4110]<= 32'hFFFFFFFF;
BRAM[4111]<= 32'hFFBAABFF;
BRAM[4112]<= 32'hFFFFFFBF;
BRAM[4113]<= 32'hFFFFFFFF;
BRAM[4114]<= 32'hFFFFFFFF;
BRAM[4115]<= 32'hF4FFFFFF;
BRAM[4116]<= 32'h00000000;
BRAM[4117]<= 32'h00000000;
BRAM[4118]<= 32'h00000000;
BRAM[4119]<= 32'hFFFFFF1B;
BRAM[4120]<= 32'hFFFFFFFF;
BRAM[4121]<= 32'hFFFFFFFF;
BRAM[4122]<= 32'hFFFFFFFF;
BRAM[4123]<= 32'hABFFFFFF;
BRAM[4124]<= 32'hFFBFFFBA;
BRAM[4125]<= 32'hFFFFFFFF;
BRAM[4126]<= 32'hFFFFFFFF;
BRAM[4127]<= 32'hFFFFFFFF;
BRAM[4128]<= 32'h0040FFFF;
BRAM[4129]<= 32'h00000000;
BRAM[4130]<= 32'h00000000;
BRAM[4131]<= 32'hFFFF0100;
BRAM[4132]<= 32'hFFFFFFFF;
BRAM[4133]<= 32'hFFFFFFFF;
BRAM[4134]<= 32'hFFFFFFFF;
BRAM[4135]<= 32'hFFFFFFFF;
BRAM[4136]<= 32'hFFBAABFF;
BRAM[4137]<= 32'hFFFFFFBF;
BRAM[4138]<= 32'hFFFFFFFF;
BRAM[4139]<= 32'hFFFFFFFF;
BRAM[4140]<= 32'hFFFFFFFF;
BRAM[4141]<= 32'h000000F4;
BRAM[4142]<= 32'h00000000;
BRAM[4143]<= 32'h1B000000;
BRAM[4144]<= 32'hFFFFFFFF;
BRAM[4145]<= 32'hFFFFFFFF;
BRAM[4146]<= 32'hFFFFFFFF;
BRAM[4147]<= 32'hFFFFFFFF;
BRAM[4148]<= 32'hABFFFFFF;
BRAM[4149]<= 32'hFFBFFFBA;
BRAM[4150]<= 32'hFFFFFFFF;
BRAM[4151]<= 32'hFFFFFFFF;
BRAM[4152]<= 32'hFFFFFFFF;
BRAM[4153]<= 32'h40FFFFFF;
BRAM[4154]<= 32'h00000000;
BRAM[4155]<= 32'h00000000;
BRAM[4156]<= 32'hFFFFBF00;
BRAM[4157]<= 32'hFFFFFFFF;
BRAM[4158]<= 32'hFFFFFFFF;
BRAM[4159]<= 32'hFFFFFFFF;
BRAM[4160]<= 32'hFFFFFFFF;
BRAM[4161]<= 32'hFFBAABFF;
BRAM[4162]<= 32'hFFFFFFBF;
BRAM[4163]<= 32'hFFFFFFFF;
BRAM[4164]<= 32'hFFFFFFFF;
BRAM[4165]<= 32'hFFFFFFFF;
BRAM[4166]<= 32'h0000E4FF;
BRAM[4167]<= 32'h00000000;
BRAM[4168]<= 32'hFF0B0000;
BRAM[4169]<= 32'hFFFFFFFF;
BRAM[4170]<= 32'hFFFFFFFF;
BRAM[4171]<= 32'hFFFFFFFF;
BRAM[4172]<= 32'hFFFFFFFF;
BRAM[4173]<= 32'hABFFFFFF;
BRAM[4174]<= 32'hFFBFFFBA;
BRAM[4175]<= 32'hFFFFFFFF;
BRAM[4176]<= 32'hFFFFFFFF;
BRAM[4177]<= 32'hFFFFFFFF;
BRAM[4178]<= 32'hFEFFFFFF;
BRAM[4179]<= 32'h00000000;
BRAM[4180]<= 32'h00000000;
BRAM[4181]<= 32'hFFFFFF7F;
BRAM[4182]<= 32'hFFFFFFFF;
BRAM[4183]<= 32'hFFFFFFFF;
BRAM[4184]<= 32'hFFFFFFFF;
BRAM[4185]<= 32'hFFFFFFFF;
BRAM[4186]<= 32'hFFBAABFF;
BRAM[4187]<= 32'hFFFFFFBF;
BRAM[4188]<= 32'hFFFFFFFF;
BRAM[4189]<= 32'hFFFFFFFF;
BRAM[4190]<= 32'hFFFFFFFF;
BRAM[4191]<= 32'h00D0FFFF;
BRAM[4192]<= 32'h00000000;
BRAM[4193]<= 32'hFFFF0700;
BRAM[4194]<= 32'hFFFFFFFF;
BRAM[4195]<= 32'hFFFFFFFF;
BRAM[4196]<= 32'hFFFFFFFF;
BRAM[4197]<= 32'hFFFFFFFF;
BRAM[4198]<= 32'hABFFFFFF;
BRAM[4199]<= 32'hFFBFFFBA;
BRAM[4200]<= 32'hFFFFFFFF;
BRAM[4201]<= 32'hFFFFFFFF;
BRAM[4202]<= 32'hFFFFFFFF;
BRAM[4203]<= 32'hFFFFFFFF;
BRAM[4204]<= 32'h000000F8;
BRAM[4205]<= 32'h2F000000;
BRAM[4206]<= 32'hFFFFFFFF;
BRAM[4207]<= 32'hFFFFFFFF;
BRAM[4208]<= 32'hFFFFFFFF;
BRAM[4209]<= 32'hFFFFFFFF;
BRAM[4210]<= 32'hFFFFFFFF;
BRAM[4211]<= 32'hFFBAABFF;
BRAM[4212]<= 32'hFFFFFFBF;
BRAM[4213]<= 32'hFFFFFFFF;
BRAM[4214]<= 32'hFFFFFFFF;
BRAM[4215]<= 32'hFFFFFFFF;
BRAM[4216]<= 32'h40FFFFFF;
BRAM[4217]<= 32'h00000000;
BRAM[4218]<= 32'hFFFFFF01;
BRAM[4219]<= 32'hFFFFFFFF;
BRAM[4220]<= 32'hFFFFFFFF;
BRAM[4221]<= 32'hFFFFFFFF;
BRAM[4222]<= 32'hFFFFFFFF;
BRAM[4223]<= 32'hABFFFFFF;
BRAM[4224]<= 32'hFFBFFFBA;
BRAM[4225]<= 32'hFFFFFFFF;
BRAM[4226]<= 32'hFFFFFFFF;
BRAM[4227]<= 32'hFFFFFFFF;
BRAM[4228]<= 32'hFFFFFFFF;
BRAM[4229]<= 32'h0000E0FF;
BRAM[4230]<= 32'hFF0B0000;
BRAM[4231]<= 32'hFFFFFFFF;
BRAM[4232]<= 32'hFFFFFFFF;
BRAM[4233]<= 32'hFFFFFFFF;
BRAM[4234]<= 32'hFFFFFFFF;
BRAM[4235]<= 32'hFFFFFFFF;
BRAM[4236]<= 32'hFFBAABFF;
BRAM[4237]<= 32'hFFFFFFBF;
BRAM[4238]<= 32'hFFFFFFFF;
BRAM[4239]<= 32'hFFFFFFFF;
BRAM[4240]<= 32'hFFFFFFFF;
BRAM[4241]<= 32'hFDFFFFFF;
BRAM[4242]<= 32'h00000000;
BRAM[4243]<= 32'hFFFFFF3F;
BRAM[4244]<= 32'hFFFFFFFF;
BRAM[4245]<= 32'hFFFFFFFF;
BRAM[4246]<= 32'hFFFFFFFF;
BRAM[4247]<= 32'hFFFFFFFF;
BRAM[4248]<= 32'hABFFFFFF;
BRAM[4249]<= 32'hFFBFFFBA;
BRAM[4250]<= 32'hFFFFFFFF;
BRAM[4251]<= 32'hFFFFFFFF;
BRAM[4252]<= 32'hFFFFFFFF;
BRAM[4253]<= 32'hFFFFFFFF;
BRAM[4254]<= 32'h0040FFFF;
BRAM[4255]<= 32'hFFFF0100;
BRAM[4256]<= 32'hFFFFFFFF;
BRAM[4257]<= 32'hFFFFFFFF;
BRAM[4258]<= 32'hFFFFFFFF;
BRAM[4259]<= 32'hFFFFFFFF;
BRAM[4260]<= 32'hFFFFFFFF;
BRAM[4261]<= 32'hFFBAABFF;
BRAM[4262]<= 32'hFFFFFFBF;
BRAM[4263]<= 32'hFFFFFFFF;
BRAM[4264]<= 32'hFFFFFFFF;
BRAM[4265]<= 32'hFFFFFFFF;
BRAM[4266]<= 32'hFFFFFFFF;
BRAM[4267]<= 32'h070000E0;
BRAM[4268]<= 32'hFFFFFFFF;
BRAM[4269]<= 32'hFFFFFFFF;
BRAM[4270]<= 32'hFFFFFFFF;
BRAM[4271]<= 32'hFFFFFFFF;
BRAM[4272]<= 32'hFFFFFFFF;
BRAM[4273]<= 32'hABFFFFFF;
BRAM[4274]<= 32'hFFBFFFBA;
BRAM[4275]<= 32'hFFFFFFFF;
BRAM[4276]<= 32'hFFFFFFFF;
BRAM[4277]<= 32'hFFFFFFFF;
BRAM[4278]<= 32'hFFFFFFFF;
BRAM[4279]<= 32'h00F8FFFF;
BRAM[4280]<= 32'hFFFF2F00;
BRAM[4281]<= 32'hFFFFFFFF;
BRAM[4282]<= 32'hFFFFFFFF;
BRAM[4283]<= 32'hFFFFFFFF;
BRAM[4284]<= 32'hFFFFFFFF;
BRAM[4285]<= 32'hFFFFFFFF;
BRAM[4286]<= 32'hFFBAABFF;
BRAM[4287]<= 32'hFFFFFFBF;
BRAM[4288]<= 32'hFFFFFFFF;
BRAM[4289]<= 32'hFFFFFFFF;
BRAM[4290]<= 32'hFFFFFFFF;
BRAM[4291]<= 32'hFFFFFFFF;
BRAM[4292]<= 32'h7F0000FE;
BRAM[4293]<= 32'hFFFFFFFF;
BRAM[4294]<= 32'hFFFFFFFF;
BRAM[4295]<= 32'hFFFFFFFF;
BRAM[4296]<= 32'hFFFFFFFF;
BRAM[4297]<= 32'hFFFFFFFF;
BRAM[4298]<= 32'hABFFFFFF;
BRAM[4299]<= 32'hFFBFFFBA;
BRAM[4300]<= 32'hFFFFFFFF;
BRAM[4301]<= 32'hFFFFFFFF;
BRAM[4302]<= 32'hFFFFFFFF;
BRAM[4303]<= 32'hFFFFFFFF;
BRAM[4304]<= 32'h80FFFFFF;
BRAM[4305]<= 32'hFFFFFF01;
BRAM[4306]<= 32'hFFFFFFFF;
BRAM[4307]<= 32'hFFFFFFFF;
BRAM[4308]<= 32'hFFFFFFFF;
BRAM[4309]<= 32'hFFFFFFFF;
BRAM[4310]<= 32'hFFFFFFFF;
BRAM[4311]<= 32'hFFBAABFF;
BRAM[4312]<= 32'hFFFFFFBF;
BRAM[4313]<= 32'hFFFFFFFF;
BRAM[4314]<= 32'hFFFFFFFF;
BRAM[4315]<= 32'hFFFFFFFF;
BRAM[4316]<= 32'hFFFFFFFF;
BRAM[4317]<= 32'hFF03D0FF;
BRAM[4318]<= 32'hFFFFFFFF;
BRAM[4319]<= 32'hFFFFFFFF;
BRAM[4320]<= 32'hFFFFFFFF;
BRAM[4321]<= 32'hFFFFFFFF;
BRAM[4322]<= 32'hFFFFFFFF;
BRAM[4323]<= 32'hABFFFFFF;
BRAM[4324]<= 32'hFFBFFFBA;
BRAM[4325]<= 32'hFFFFFFFF;
BRAM[4326]<= 32'hFFFFFFFF;
BRAM[4327]<= 32'hFFFFFFFF;
BRAM[4328]<= 32'hFFFFFFFF;
BRAM[4329]<= 32'hF0FFFFFF;
BRAM[4330]<= 32'hFFFFFF0F;
BRAM[4331]<= 32'hFFFFFFFF;
BRAM[4332]<= 32'hFFFFFFFF;
BRAM[4333]<= 32'hFFFFFFFF;
BRAM[4334]<= 32'hFFFFFFFF;
BRAM[4335]<= 32'hFFFFFFFF;
BRAM[4336]<= 32'hEFBAABFF;
BRAM[4337]<= 32'hFFFFFFBF;
BRAM[4338]<= 32'hFFFFFFFF;
BRAM[4339]<= 32'hFFFFFFFF;
BRAM[4340]<= 32'hFFFFFFFF;
BRAM[4341]<= 32'hFFFFFFFF;
BRAM[4342]<= 32'hFF1FF8FF;
BRAM[4343]<= 32'hFFFFFFFF;
BRAM[4344]<= 32'hFFFFFFFF;
BRAM[4345]<= 32'hFFFFFFFF;
BRAM[4346]<= 32'hFFFFFFFF;
BRAM[4347]<= 32'hFFFFFFFF;
BRAM[4348]<= 32'hFFFFFFFF;
BRAM[4349]<= 32'hFFFFFFFF;
BRAM[4350]<= 32'hFFFFFFFF;
BRAM[4351]<= 32'hFFFFFFFF;
BRAM[4352]<= 32'hFFFFFFFF;
BRAM[4353]<= 32'hFFFFFFFF;
BRAM[4354]<= 32'hFCFFFFFF;
BRAM[4355]<= 32'hFFFFFF3F;
BRAM[4356]<= 32'hFFFFFFFF;
BRAM[4357]<= 32'hFFFFFFFF;
BRAM[4358]<= 32'hFFFFFFFF;
BRAM[4359]<= 32'hFFFFFFFF;
BRAM[4360]<= 32'hFFFFFFFF;
BRAM[4361]<= 32'hFFFFFFFF;
BRAM[4362]<= 32'hFFFFFFFF;
BRAM[4363]<= 32'hFFFFFFFF;
BRAM[4364]<= 32'hFFFFFFFF;
BRAM[4365]<= 32'hFFFFFFFF;
BRAM[4366]<= 32'hFFFFFFFF;
BRAM[4367]<= 32'hFFFFFFFF;
BRAM[4368]<= 32'hFFFFFFFF;
BRAM[4369]<= 32'hFFFFFFFF;
BRAM[4370]<= 32'hFFFFFFFF;
BRAM[4371]<= 32'hFFFFFFFF;
BRAM[4372]<= 32'hFFFFFFFF;
BRAM[4373]<= 32'hFFFFFFFF;
BRAM[4374]<= 32'hFFFFFFFF;
BRAM[4375]<= 32'hFFFFFFFF;
BRAM[4376]<= 32'hFFFFFFFF;
BRAM[4377]<= 32'hFFFFFFFF;
BRAM[4378]<= 32'hFFFFFFFF;
BRAM[4379]<= 32'hFFFFFFFF;
BRAM[4380]<= 32'hFFFFFFFF;
BRAM[4381]<= 32'hFFFFFFFF;
BRAM[4382]<= 32'hFFFFFFFF;
BRAM[4383]<= 32'hFFFFFFFF;
BRAM[4384]<= 32'hFFFFFFFF;
BRAM[4385]<= 32'hFFFFFFFF;
BRAM[4386]<= 32'h00000000;
BRAM[4387]<= 32'h00000000;
BRAM[4388]<= 32'h80110000;
BRAM[4389]<= 32'h00000000;
BRAM[4390]<= 32'h00000000;
BRAM[4391]<= 32'h00000000;
BRAM[4392]<= 32'h00000000;
BRAM[4393]<= 32'hC0070000;
BRAM[4394]<= 32'h8003FC7F;
BRAM[4395]<= 32'h80319C33;
BRAM[4396]<= 32'hE600FE3F;
BRAM[4397]<= 32'hFE7E8001;
BRAM[4398]<= 32'h3F0E060E;
BRAM[4399]<= 32'h7003060E;
BRAM[4400]<= 32'hFE3FC001;
BRAM[4401]<= 32'h0C60F03F;
BRAM[4402]<= 32'hFE7F8001;
BRAM[4403]<= 32'hC061FC73;
BRAM[4404]<= 32'hFC3FF63F;
BRAM[4405]<= 32'h363FC666;
BRAM[4406]<= 32'h363FB03F;
BRAM[4407]<= 32'hC0007773;
BRAM[4408]<= 32'h3CF81736;
BRAM[4409]<= 32'hFC7FE44F;
BRAM[4410]<= 32'hFC7F0660;
BRAM[4411]<= 32'h6030FCFF;
BRAM[4412]<= 32'hC6668E71;
BRAM[4413]<= 32'h3031B673;
BRAM[4414]<= 32'h7733B67B;
BRAM[4415]<= 32'h3806FE3F;
BRAM[4416]<= 32'h8C430EE0;
BRAM[4417]<= 32'h0660FC7F;
BRAM[4418]<= 32'hC0718061;
BRAM[4419]<= 32'h86316430;
BRAM[4420]<= 32'hB6603E66;
BRAM[4421]<= 32'h9660303B;
BRAM[4422]<= 32'hFE3F7633;
BRAM[4423]<= 32'hF83FFC0F;
BRAM[4424]<= 32'h00010C61;
BRAM[4425]<= 32'h80E1001F;
BRAM[4426]<= 32'h6438C071;
BRAM[4427]<= 32'h7C668E71;
BRAM[4428]<= 32'hBF7F3640;
BRAM[4429]<= 32'h76333600;
BRAM[4430]<= 32'h3A0EC000;
BRAM[4431]<= 32'h8C638003;
BRAM[4432]<= 32'hF81F8001;
BRAM[4433]<= 32'hFC7F8001;
BRAM[4434]<= 32'hFE7F683E;
BRAM[4435]<= 32'hB67FFE7E;
BRAM[4436]<= 32'hB63F3600;
BRAM[4437]<= 32'hC0007633;
BRAM[4438]<= 32'h00033A06;
BRAM[4439]<= 32'h8003E44F;
BRAM[4440]<= 32'h8001F000;
BRAM[4441]<= 32'h7836C061;
BRAM[4442]<= 32'h820C8E71;
BRAM[4443]<= 32'h360CB671;
BRAM[4444]<= 32'h7633B631;
BRAM[4445]<= 32'hF927C001;
BRAM[4446]<= 32'h0C630003;
BRAM[4447]<= 32'hC001C007;
BRAM[4448]<= 32'hFE7FFC3F;
BRAM[4449]<= 32'h86313036;
BRAM[4450]<= 32'hB671102C;
BRAM[4451]<= 32'hB631B63F;
BRAM[4452]<= 32'hE0036633;
BRAM[4453]<= 32'hFC7F0E3C;
BRAM[4454]<= 32'hE00E2C61;
BRAM[4455]<= 32'h8001FE7F;
BRAM[4456]<= 32'h30360000;
BRAM[4457]<= 32'hFE6EFE77;
BRAM[4458]<= 32'h360CB677;
BRAM[4459]<= 32'h6633B637;
BRAM[4460]<= 32'h2E3E7007;
BRAM[4461]<= 32'hA4630003;
BRAM[4462]<= 32'h8001701C;
BRAM[4463]<= 32'hFE5F8001;
BRAM[4464]<= 32'hF83F3636;
BRAM[4465]<= 32'h3676C66C;
BRAM[4466]<= 32'h3636362F;
BRAM[4467]<= 32'h38066E3B;
BRAM[4468]<= 32'h0003CE18;
BRAM[4469]<= 32'h3018F45F;
BRAM[4470]<= 32'h80018001;
BRAM[4471]<= 32'h7E368001;
BRAM[4472]<= 32'hC66C8001;
BRAM[4473]<= 32'hB62D8670;
BRAM[4474]<= 32'h6003C630;
BRAM[4475]<= 32'hC618180E;
BRAM[4476]<= 32'h0C400003;
BRAM[4477]<= 32'h80013838;
BRAM[4478]<= 32'h9C398001;
BRAM[4479]<= 32'h86015E6E;
BRAM[4480]<= 32'h8671C66C;
BRAM[4481]<= 32'h8631B66D;
BRAM[4482]<= 32'h1C1C7003;
BRAM[4483]<= 32'hFCFFFC0F;
BRAM[4484]<= 32'h1C70FEFF;
BRAM[4485]<= 32'hFE7F8007;
BRAM[4486]<= 32'hCC608E71;
BRAM[4487]<= 32'hFE7EFE01;
BRAM[4488]<= 32'hE66D9E7F;
BRAM[4489]<= 32'hFF7F9E7F;
BRAM[4490]<= 32'h3F3F0E38;
BRAM[4491]<= 32'h00000000;
BRAM[4492]<= 32'h00000000;
BRAM[4493]<= 32'h00000000;
BRAM[4494]<= 32'h00008000;
BRAM[4495]<= 32'h00000000;
BRAM[4496]<= 32'h00000000;
BRAM[4497]<= 32'h00000000;
BRAM[4498]<= 32'h00000000;
BRAM[4499]<= 32'h00000000;
BRAM[4500]<= 32'h00000000;
BRAM[4501]<= 32'h00000000;
BRAM[4502]<= 32'h00000000;
BRAM[4503]<= 32'h00000000;
BRAM[4504]<= 32'h00000000;
BRAM[4505]<= 32'h00000000;
BRAM[4506]<= 32'h00000000;
BRAM[4507]<= 32'h00000000;
BRAM[4508]<= 32'h00000000;
BRAM[4509]<= 32'h00000000;
BRAM[4510]<= 32'h00000000;
BRAM[4511]<= 32'h00000000;
BRAM[4512]<= 32'h00000000;
BRAM[4513]<= 32'h00000000;
BRAM[4514]<= 32'h00000000;
BRAM[4515]<= 32'h00000000;
BRAM[4516]<= 32'h00000000;
BRAM[4517]<= 32'h00000000;
BRAM[4518]<= 32'h00000000;
BRAM[4519]<= 32'h00000000;
BRAM[4520]<= 32'h00000000;
BRAM[4521]<= 32'h0887203E;
BRAM[4522]<= 32'hC1034060;
BRAM[4523]<= 32'h7C8080E0;
BRAM[4524]<= 32'h70800F1E;
BRAM[4525]<= 32'hF0E10178;
BRAM[4526]<= 32'hE3838741;
BRAM[4527]<= 32'hE1F1E3F8;
BRAM[4528]<= 32'h206041F0;
BRAM[4529]<= 32'hE0600C82;
BRAM[4530]<= 32'h80100204;
BRAM[4531]<= 32'h0820C080;
BRAM[4532]<= 32'h02C02000;
BRAM[4533]<= 32'h84611803;
BRAM[4534]<= 32'h40400042;
BRAM[4535]<= 32'h61184140;
BRAM[4536]<= 32'h0A822040;
BRAM[4537]<= 32'h040CA060;
BRAM[4538]<= 32'hC0808010;
BRAM[4539]<= 32'h20000840;
BRAM[4540]<= 32'h08020480;
BRAM[4541]<= 32'h00428452;
BRAM[4542]<= 32'h42404040;
BRAM[4543]<= 32'h3F405108;
BRAM[4544]<= 32'h10610B82;
BRAM[4545]<= 32'h80080408;
BRAM[4546]<= 32'h0F407880;
BRAM[4547]<= 32'h04802080;
BRAM[4548]<= 32'h875C0802;
BRAM[4549]<= 32'h4040E0C3;
BRAM[4550]<= 32'h49084240;
BRAM[4551]<= 32'h09822040;
BRAM[4552]<= 32'h040CF0E1;
BRAM[4553]<= 32'hC0808010;
BRAM[4554]<= 32'h20000841;
BRAM[4555]<= 32'h08020480;
BRAM[4556]<= 32'h00028748;
BRAM[4557]<= 32'h42404040;
BRAM[4558]<= 32'h20604508;
BRAM[4559]<= 32'h08E20882;
BRAM[4560]<= 32'h80100204;
BRAM[4561]<= 32'h0821C080;
BRAM[4562]<= 32'h02C02000;
BRAM[4563]<= 32'h84401803;
BRAM[4564]<= 32'h40400002;
BRAM[4565]<= 32'h47184140;
BRAM[4566]<= 32'h0887203E;
BRAM[4567]<= 32'hC1030842;
BRAM[4568]<= 32'h7CF8F8E0;
BRAM[4569]<= 32'h70800F1F;
BRAM[4570]<= 32'hF0E1017C;
BRAM[4571]<= 32'hE0038440;
BRAM[4572]<= 32'hE141E040;
BRAM[4573]<= 32'h000043F0;
BRAM[4574]<= 32'h00004798;
BRAM[4575]<= 32'h20000000;
BRAM[4576]<= 32'h0000001C;
BRAM[4577]<= 32'h0000008C;
BRAM[4578]<= 32'h000047B4;
BRAM[4579]<= 32'h2000001C;
BRAM[4580]<= 32'h0000A064;
BRAM[4581]<= 32'h000000A8;
BRAM[4582]<= 32'h00000000;
BRAM[4583]<= 32'h00000000;
BRAM[4584]<= 32'h00000000;
BRAM[4585]<= 32'h00000000;
BRAM[4586]<= 32'h00000000;
BRAM[4587]<= 32'h00000000;
BRAM[4588]<= 32'h02FAF080;
end